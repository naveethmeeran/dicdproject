magic
tech scmos
timestamp 1509121979
<< ab >>
rect 16 235 56 379
rect 58 235 185 379
rect 193 235 320 379
rect 322 235 362 379
rect 363 235 490 379
rect 492 235 572 379
rect 574 235 701 379
rect 16 163 400 235
rect 14 155 400 163
rect 11 91 400 155
rect 413 91 701 235
rect 16 19 56 91
rect 57 19 399 91
rect 412 19 700 91
<< nwell >>
rect 11 339 705 384
rect 11 195 705 275
rect 11 51 705 131
<< pwell >>
rect 11 275 705 339
rect 11 131 705 195
rect 11 14 705 51
<< poly >>
rect 25 373 27 377
rect 35 373 37 377
rect 45 373 47 377
rect 65 373 67 377
rect 75 373 77 377
rect 85 373 87 377
rect 106 373 108 377
rect 116 373 118 377
rect 126 373 128 377
rect 25 350 27 354
rect 21 348 27 350
rect 21 346 23 348
rect 25 346 27 348
rect 21 344 27 346
rect 25 333 27 344
rect 35 342 37 354
rect 65 350 67 354
rect 61 348 67 350
rect 61 346 63 348
rect 65 346 67 348
rect 45 342 47 345
rect 61 344 67 346
rect 31 340 37 342
rect 31 338 33 340
rect 35 338 37 340
rect 31 336 37 338
rect 41 340 47 342
rect 41 338 43 340
rect 45 338 47 340
rect 41 336 47 338
rect 32 333 34 336
rect 45 333 47 336
rect 65 333 67 344
rect 75 342 77 354
rect 144 370 146 375
rect 151 370 153 375
rect 174 373 176 377
rect 202 373 204 377
rect 161 361 163 366
rect 225 370 227 375
rect 232 370 234 375
rect 250 373 252 377
rect 260 373 262 377
rect 270 373 272 377
rect 291 373 293 377
rect 301 373 303 377
rect 311 373 313 377
rect 331 373 333 377
rect 341 373 343 377
rect 351 373 353 377
rect 372 373 374 377
rect 215 361 217 366
rect 161 345 163 348
rect 85 342 87 345
rect 106 342 108 345
rect 116 342 118 345
rect 126 342 128 345
rect 144 342 146 345
rect 151 342 153 345
rect 161 343 170 345
rect 71 340 77 342
rect 71 338 73 340
rect 75 338 77 340
rect 71 336 77 338
rect 81 340 87 342
rect 81 338 83 340
rect 85 338 87 340
rect 81 336 87 338
rect 104 340 110 342
rect 104 338 106 340
rect 108 338 110 340
rect 104 336 110 338
rect 114 340 120 342
rect 114 338 116 340
rect 118 338 120 340
rect 114 336 120 338
rect 124 340 146 342
rect 124 338 126 340
rect 128 338 133 340
rect 135 338 146 340
rect 124 336 146 338
rect 150 340 156 342
rect 150 338 152 340
rect 154 338 156 340
rect 150 336 156 338
rect 72 333 74 336
rect 85 333 87 336
rect 25 315 27 320
rect 32 315 34 320
rect 45 314 47 319
rect 65 315 67 320
rect 72 315 74 320
rect 106 327 108 336
rect 117 333 119 336
rect 124 333 126 336
rect 144 333 146 336
rect 154 333 156 336
rect 164 341 166 343
rect 168 341 170 343
rect 164 339 170 341
rect 85 314 87 319
rect 164 326 166 339
rect 174 335 176 348
rect 170 333 176 335
rect 170 331 172 333
rect 174 331 176 333
rect 170 329 176 331
rect 174 326 176 329
rect 202 335 204 348
rect 215 345 217 348
rect 208 343 217 345
rect 208 341 210 343
rect 212 341 214 343
rect 225 342 227 345
rect 232 342 234 345
rect 250 342 252 345
rect 260 342 262 345
rect 270 342 272 345
rect 291 342 293 345
rect 301 342 303 354
rect 311 350 313 354
rect 311 348 317 350
rect 311 346 313 348
rect 315 346 317 348
rect 311 344 317 346
rect 208 339 214 341
rect 202 333 208 335
rect 202 331 204 333
rect 206 331 208 333
rect 202 329 208 331
rect 202 326 204 329
rect 212 326 214 339
rect 222 340 228 342
rect 222 338 224 340
rect 226 338 228 340
rect 222 336 228 338
rect 232 340 254 342
rect 232 338 243 340
rect 245 338 250 340
rect 252 338 254 340
rect 232 336 254 338
rect 258 340 264 342
rect 258 338 260 340
rect 262 338 264 340
rect 258 336 264 338
rect 268 340 274 342
rect 268 338 270 340
rect 272 338 274 340
rect 268 336 274 338
rect 291 340 297 342
rect 291 338 293 340
rect 295 338 297 340
rect 291 336 297 338
rect 301 340 307 342
rect 301 338 303 340
rect 305 338 307 340
rect 301 336 307 338
rect 222 333 224 336
rect 232 333 234 336
rect 252 333 254 336
rect 259 333 261 336
rect 144 314 146 319
rect 154 314 156 319
rect 106 309 108 313
rect 117 309 119 313
rect 124 309 126 313
rect 164 311 166 316
rect 174 309 176 313
rect 202 309 204 313
rect 212 311 214 316
rect 222 314 224 319
rect 232 314 234 319
rect 270 327 272 336
rect 291 333 293 336
rect 304 333 306 336
rect 311 333 313 344
rect 331 342 333 345
rect 341 342 343 354
rect 351 350 353 354
rect 351 348 357 350
rect 395 370 397 375
rect 402 370 404 375
rect 420 373 422 377
rect 430 373 432 377
rect 440 373 442 377
rect 461 373 463 377
rect 471 373 473 377
rect 481 373 483 377
rect 501 373 503 377
rect 511 373 513 377
rect 521 373 523 377
rect 541 373 543 377
rect 551 373 553 377
rect 561 373 563 377
rect 581 373 583 377
rect 591 373 593 377
rect 601 373 603 377
rect 622 373 624 377
rect 632 373 634 377
rect 642 373 644 377
rect 385 361 387 366
rect 351 346 353 348
rect 355 346 357 348
rect 351 344 357 346
rect 331 340 337 342
rect 331 338 333 340
rect 335 338 337 340
rect 331 336 337 338
rect 341 340 347 342
rect 341 338 343 340
rect 345 338 347 340
rect 341 336 347 338
rect 331 333 333 336
rect 344 333 346 336
rect 351 333 353 344
rect 372 335 374 348
rect 385 345 387 348
rect 378 343 387 345
rect 378 341 380 343
rect 382 341 384 343
rect 395 342 397 345
rect 402 342 404 345
rect 420 342 422 345
rect 430 342 432 345
rect 440 342 442 345
rect 461 342 463 345
rect 471 342 473 354
rect 481 350 483 354
rect 481 348 487 350
rect 481 346 483 348
rect 485 346 487 348
rect 481 344 487 346
rect 378 339 384 341
rect 372 333 378 335
rect 291 314 293 319
rect 304 315 306 320
rect 311 315 313 320
rect 372 331 374 333
rect 376 331 378 333
rect 372 329 378 331
rect 372 326 374 329
rect 382 326 384 339
rect 392 340 398 342
rect 392 338 394 340
rect 396 338 398 340
rect 392 336 398 338
rect 402 340 424 342
rect 402 338 413 340
rect 415 338 420 340
rect 422 338 424 340
rect 402 336 424 338
rect 428 340 434 342
rect 428 338 430 340
rect 432 338 434 340
rect 428 336 434 338
rect 438 340 444 342
rect 438 338 440 340
rect 442 338 444 340
rect 438 336 444 338
rect 461 340 467 342
rect 461 338 463 340
rect 465 338 467 340
rect 461 336 467 338
rect 471 340 477 342
rect 471 338 473 340
rect 475 338 477 340
rect 471 336 477 338
rect 392 333 394 336
rect 402 333 404 336
rect 422 333 424 336
rect 429 333 431 336
rect 331 314 333 319
rect 344 315 346 320
rect 351 315 353 320
rect 252 309 254 313
rect 259 309 261 313
rect 270 309 272 313
rect 372 309 374 313
rect 382 311 384 316
rect 392 314 394 319
rect 402 314 404 319
rect 440 327 442 336
rect 461 333 463 336
rect 474 333 476 336
rect 481 333 483 344
rect 501 342 503 345
rect 511 342 513 354
rect 521 350 523 354
rect 541 350 543 354
rect 521 348 527 350
rect 521 346 523 348
rect 525 346 527 348
rect 521 344 527 346
rect 537 348 543 350
rect 537 346 539 348
rect 541 346 543 348
rect 537 344 543 346
rect 501 340 507 342
rect 501 338 503 340
rect 505 338 507 340
rect 501 336 507 338
rect 511 340 517 342
rect 511 338 513 340
rect 515 338 517 340
rect 511 336 517 338
rect 501 333 503 336
rect 514 333 516 336
rect 521 333 523 344
rect 541 333 543 344
rect 551 342 553 354
rect 581 350 583 354
rect 577 348 583 350
rect 577 346 579 348
rect 581 346 583 348
rect 561 342 563 345
rect 577 344 583 346
rect 547 340 553 342
rect 547 338 549 340
rect 551 338 553 340
rect 547 336 553 338
rect 557 340 563 342
rect 557 338 559 340
rect 561 338 563 340
rect 557 336 563 338
rect 548 333 550 336
rect 561 333 563 336
rect 581 333 583 344
rect 591 342 593 354
rect 660 370 662 375
rect 667 370 669 375
rect 690 373 692 377
rect 677 361 679 366
rect 677 345 679 348
rect 601 342 603 345
rect 622 342 624 345
rect 632 342 634 345
rect 642 342 644 345
rect 660 342 662 345
rect 667 342 669 345
rect 677 343 686 345
rect 587 340 593 342
rect 587 338 589 340
rect 591 338 593 340
rect 587 336 593 338
rect 597 340 603 342
rect 597 338 599 340
rect 601 338 603 340
rect 597 336 603 338
rect 620 340 626 342
rect 620 338 622 340
rect 624 338 626 340
rect 620 336 626 338
rect 630 340 636 342
rect 630 338 632 340
rect 634 338 636 340
rect 630 336 636 338
rect 640 340 662 342
rect 640 338 642 340
rect 644 338 649 340
rect 651 338 662 340
rect 640 336 662 338
rect 666 340 672 342
rect 666 338 668 340
rect 670 338 672 340
rect 666 336 672 338
rect 588 333 590 336
rect 601 333 603 336
rect 461 314 463 319
rect 474 315 476 320
rect 481 315 483 320
rect 501 314 503 319
rect 514 315 516 320
rect 521 315 523 320
rect 541 315 543 320
rect 548 315 550 320
rect 422 309 424 313
rect 429 309 431 313
rect 440 309 442 313
rect 561 314 563 319
rect 581 315 583 320
rect 588 315 590 320
rect 622 327 624 336
rect 633 333 635 336
rect 640 333 642 336
rect 660 333 662 336
rect 670 333 672 336
rect 680 341 682 343
rect 684 341 686 343
rect 680 339 686 341
rect 601 314 603 319
rect 680 326 682 339
rect 690 335 692 348
rect 686 333 692 335
rect 686 331 688 333
rect 690 331 692 333
rect 686 329 692 331
rect 690 326 692 329
rect 660 314 662 319
rect 670 314 672 319
rect 622 309 624 313
rect 633 309 635 313
rect 640 309 642 313
rect 680 311 682 316
rect 690 309 692 313
rect 106 301 108 305
rect 117 301 119 305
rect 124 301 126 305
rect 25 294 27 299
rect 32 294 34 299
rect 45 295 47 300
rect 65 294 67 299
rect 72 294 74 299
rect 85 295 87 300
rect 25 270 27 281
rect 32 278 34 281
rect 45 278 47 281
rect 31 276 37 278
rect 31 274 33 276
rect 35 274 37 276
rect 31 272 37 274
rect 41 276 47 278
rect 41 274 43 276
rect 45 274 47 276
rect 41 272 47 274
rect 21 268 27 270
rect 21 266 23 268
rect 25 266 27 268
rect 21 264 27 266
rect 25 260 27 264
rect 35 260 37 272
rect 45 269 47 272
rect 65 270 67 281
rect 72 278 74 281
rect 85 278 87 281
rect 106 278 108 287
rect 144 295 146 300
rect 154 295 156 300
rect 164 298 166 303
rect 174 301 176 305
rect 202 301 204 305
rect 212 298 214 303
rect 252 301 254 305
rect 259 301 261 305
rect 270 301 272 305
rect 222 295 224 300
rect 232 295 234 300
rect 117 278 119 281
rect 124 278 126 281
rect 144 278 146 281
rect 154 278 156 281
rect 71 276 77 278
rect 71 274 73 276
rect 75 274 77 276
rect 71 272 77 274
rect 81 276 87 278
rect 81 274 83 276
rect 85 274 87 276
rect 81 272 87 274
rect 104 276 110 278
rect 104 274 106 276
rect 108 274 110 276
rect 104 272 110 274
rect 114 276 120 278
rect 114 274 116 276
rect 118 274 120 276
rect 114 272 120 274
rect 124 276 146 278
rect 124 274 126 276
rect 128 274 133 276
rect 135 274 146 276
rect 124 272 146 274
rect 150 276 156 278
rect 150 274 152 276
rect 154 274 156 276
rect 150 272 156 274
rect 164 275 166 288
rect 174 285 176 288
rect 170 283 176 285
rect 170 281 172 283
rect 174 281 176 283
rect 170 279 176 281
rect 164 273 170 275
rect 61 268 67 270
rect 61 266 63 268
rect 65 266 67 268
rect 61 264 67 266
rect 65 260 67 264
rect 75 260 77 272
rect 85 269 87 272
rect 106 269 108 272
rect 116 269 118 272
rect 126 269 128 272
rect 144 269 146 272
rect 151 269 153 272
rect 164 271 166 273
rect 168 271 170 273
rect 161 269 170 271
rect 161 266 163 269
rect 174 266 176 279
rect 202 285 204 288
rect 202 283 208 285
rect 202 281 204 283
rect 206 281 208 283
rect 202 279 208 281
rect 202 266 204 279
rect 212 275 214 288
rect 372 301 374 305
rect 291 295 293 300
rect 208 273 214 275
rect 208 271 210 273
rect 212 271 214 273
rect 222 278 224 281
rect 232 278 234 281
rect 252 278 254 281
rect 259 278 261 281
rect 270 278 272 287
rect 304 294 306 299
rect 311 294 313 299
rect 331 295 333 300
rect 344 294 346 299
rect 351 294 353 299
rect 382 298 384 303
rect 422 301 424 305
rect 429 301 431 305
rect 440 301 442 305
rect 392 295 394 300
rect 402 295 404 300
rect 372 285 374 288
rect 372 283 378 285
rect 372 281 374 283
rect 376 281 378 283
rect 291 278 293 281
rect 304 278 306 281
rect 222 276 228 278
rect 222 274 224 276
rect 226 274 228 276
rect 222 272 228 274
rect 232 276 254 278
rect 232 274 243 276
rect 245 274 250 276
rect 252 274 254 276
rect 232 272 254 274
rect 258 276 264 278
rect 258 274 260 276
rect 262 274 264 276
rect 258 272 264 274
rect 268 276 274 278
rect 268 274 270 276
rect 272 274 274 276
rect 268 272 274 274
rect 291 276 297 278
rect 291 274 293 276
rect 295 274 297 276
rect 291 272 297 274
rect 301 276 307 278
rect 301 274 303 276
rect 305 274 307 276
rect 301 272 307 274
rect 208 269 217 271
rect 225 269 227 272
rect 232 269 234 272
rect 250 269 252 272
rect 260 269 262 272
rect 270 269 272 272
rect 291 269 293 272
rect 215 266 217 269
rect 161 248 163 253
rect 25 237 27 241
rect 35 237 37 241
rect 45 237 47 241
rect 65 237 67 241
rect 75 237 77 241
rect 85 237 87 241
rect 106 237 108 241
rect 116 237 118 241
rect 126 237 128 241
rect 144 239 146 244
rect 151 239 153 244
rect 215 248 217 253
rect 174 237 176 241
rect 202 237 204 241
rect 225 239 227 244
rect 232 239 234 244
rect 301 260 303 272
rect 311 270 313 281
rect 331 278 333 281
rect 344 278 346 281
rect 331 276 337 278
rect 331 274 333 276
rect 335 274 337 276
rect 331 272 337 274
rect 341 276 347 278
rect 341 274 343 276
rect 345 274 347 276
rect 341 272 347 274
rect 311 268 317 270
rect 331 269 333 272
rect 311 266 313 268
rect 315 266 317 268
rect 311 264 317 266
rect 311 260 313 264
rect 341 260 343 272
rect 351 270 353 281
rect 372 279 378 281
rect 351 268 357 270
rect 351 266 353 268
rect 355 266 357 268
rect 372 266 374 279
rect 382 275 384 288
rect 461 295 463 300
rect 378 273 384 275
rect 378 271 380 273
rect 382 271 384 273
rect 392 278 394 281
rect 402 278 404 281
rect 422 278 424 281
rect 429 278 431 281
rect 440 278 442 287
rect 474 294 476 299
rect 481 294 483 299
rect 501 295 503 300
rect 622 301 624 305
rect 633 301 635 305
rect 640 301 642 305
rect 514 294 516 299
rect 521 294 523 299
rect 541 294 543 299
rect 548 294 550 299
rect 561 295 563 300
rect 581 294 583 299
rect 588 294 590 299
rect 601 295 603 300
rect 461 278 463 281
rect 474 278 476 281
rect 392 276 398 278
rect 392 274 394 276
rect 396 274 398 276
rect 392 272 398 274
rect 402 276 424 278
rect 402 274 413 276
rect 415 274 420 276
rect 422 274 424 276
rect 402 272 424 274
rect 428 276 434 278
rect 428 274 430 276
rect 432 274 434 276
rect 428 272 434 274
rect 438 276 444 278
rect 438 274 440 276
rect 442 274 444 276
rect 438 272 444 274
rect 461 276 467 278
rect 461 274 463 276
rect 465 274 467 276
rect 461 272 467 274
rect 471 276 477 278
rect 471 274 473 276
rect 475 274 477 276
rect 471 272 477 274
rect 378 269 387 271
rect 395 269 397 272
rect 402 269 404 272
rect 420 269 422 272
rect 430 269 432 272
rect 440 269 442 272
rect 461 269 463 272
rect 385 266 387 269
rect 351 264 357 266
rect 351 260 353 264
rect 385 248 387 253
rect 250 237 252 241
rect 260 237 262 241
rect 270 237 272 241
rect 291 237 293 241
rect 301 237 303 241
rect 311 237 313 241
rect 331 237 333 241
rect 341 237 343 241
rect 351 237 353 241
rect 372 237 374 241
rect 395 239 397 244
rect 402 239 404 244
rect 471 260 473 272
rect 481 270 483 281
rect 501 278 503 281
rect 514 278 516 281
rect 501 276 507 278
rect 501 274 503 276
rect 505 274 507 276
rect 501 272 507 274
rect 511 276 517 278
rect 511 274 513 276
rect 515 274 517 276
rect 511 272 517 274
rect 481 268 487 270
rect 501 269 503 272
rect 481 266 483 268
rect 485 266 487 268
rect 481 264 487 266
rect 481 260 483 264
rect 511 260 513 272
rect 521 270 523 281
rect 541 270 543 281
rect 548 278 550 281
rect 561 278 563 281
rect 547 276 553 278
rect 547 274 549 276
rect 551 274 553 276
rect 547 272 553 274
rect 557 276 563 278
rect 557 274 559 276
rect 561 274 563 276
rect 557 272 563 274
rect 521 268 527 270
rect 521 266 523 268
rect 525 266 527 268
rect 521 264 527 266
rect 537 268 543 270
rect 537 266 539 268
rect 541 266 543 268
rect 537 264 543 266
rect 521 260 523 264
rect 541 260 543 264
rect 551 260 553 272
rect 561 269 563 272
rect 581 270 583 281
rect 588 278 590 281
rect 601 278 603 281
rect 622 278 624 287
rect 660 295 662 300
rect 670 295 672 300
rect 680 298 682 303
rect 690 301 692 305
rect 633 278 635 281
rect 640 278 642 281
rect 660 278 662 281
rect 670 278 672 281
rect 587 276 593 278
rect 587 274 589 276
rect 591 274 593 276
rect 587 272 593 274
rect 597 276 603 278
rect 597 274 599 276
rect 601 274 603 276
rect 597 272 603 274
rect 620 276 626 278
rect 620 274 622 276
rect 624 274 626 276
rect 620 272 626 274
rect 630 276 636 278
rect 630 274 632 276
rect 634 274 636 276
rect 630 272 636 274
rect 640 276 662 278
rect 640 274 642 276
rect 644 274 649 276
rect 651 274 662 276
rect 640 272 662 274
rect 666 276 672 278
rect 666 274 668 276
rect 670 274 672 276
rect 666 272 672 274
rect 680 275 682 288
rect 690 285 692 288
rect 686 283 692 285
rect 686 281 688 283
rect 690 281 692 283
rect 686 279 692 281
rect 680 273 686 275
rect 577 268 583 270
rect 577 266 579 268
rect 581 266 583 268
rect 577 264 583 266
rect 581 260 583 264
rect 591 260 593 272
rect 601 269 603 272
rect 622 269 624 272
rect 632 269 634 272
rect 642 269 644 272
rect 660 269 662 272
rect 667 269 669 272
rect 680 271 682 273
rect 684 271 686 273
rect 677 269 686 271
rect 677 266 679 269
rect 690 266 692 279
rect 677 248 679 253
rect 420 237 422 241
rect 430 237 432 241
rect 440 237 442 241
rect 461 237 463 241
rect 471 237 473 241
rect 481 237 483 241
rect 501 237 503 241
rect 511 237 513 241
rect 521 237 523 241
rect 541 237 543 241
rect 551 237 553 241
rect 561 237 563 241
rect 581 237 583 241
rect 591 237 593 241
rect 601 237 603 241
rect 622 237 624 241
rect 632 237 634 241
rect 642 237 644 241
rect 660 239 662 244
rect 667 239 669 244
rect 690 237 692 241
rect 25 229 27 233
rect 38 229 40 233
rect 45 229 47 233
rect 66 229 68 233
rect 76 229 78 233
rect 86 229 88 233
rect 104 226 106 231
rect 111 226 113 231
rect 134 229 136 233
rect 167 229 169 233
rect 177 229 179 233
rect 187 229 189 233
rect 121 217 123 222
rect 121 201 123 204
rect 25 198 27 201
rect 38 198 40 201
rect 45 198 47 201
rect 66 198 68 201
rect 76 198 78 201
rect 86 198 88 201
rect 104 198 106 201
rect 111 198 113 201
rect 121 199 130 201
rect 25 196 31 198
rect 25 194 27 196
rect 29 194 31 196
rect 25 192 31 194
rect 35 196 41 198
rect 35 194 37 196
rect 39 194 41 196
rect 35 192 41 194
rect 45 196 54 198
rect 45 194 50 196
rect 52 194 54 196
rect 45 192 54 194
rect 64 196 70 198
rect 64 194 66 196
rect 68 194 70 196
rect 64 192 70 194
rect 74 196 80 198
rect 74 194 76 196
rect 78 194 80 196
rect 74 192 80 194
rect 84 196 106 198
rect 84 194 86 196
rect 88 194 93 196
rect 95 194 106 196
rect 84 192 106 194
rect 110 196 116 198
rect 110 194 112 196
rect 114 194 116 196
rect 110 192 116 194
rect 25 189 27 192
rect 35 184 37 192
rect 45 186 47 192
rect 66 183 68 192
rect 77 189 79 192
rect 84 189 86 192
rect 104 189 106 192
rect 114 189 116 192
rect 124 197 126 199
rect 128 197 130 199
rect 124 195 130 197
rect 25 170 27 175
rect 35 171 37 176
rect 45 174 47 178
rect 124 182 126 195
rect 134 191 136 204
rect 205 226 207 231
rect 212 226 214 231
rect 235 229 237 233
rect 269 229 271 233
rect 279 229 281 233
rect 289 229 291 233
rect 222 217 224 222
rect 222 201 224 204
rect 167 198 169 201
rect 177 198 179 201
rect 187 198 189 201
rect 205 198 207 201
rect 212 198 214 201
rect 222 199 231 201
rect 165 196 171 198
rect 165 194 167 196
rect 169 194 171 196
rect 165 192 171 194
rect 175 196 181 198
rect 175 194 177 196
rect 179 194 181 196
rect 175 192 181 194
rect 185 196 207 198
rect 185 194 187 196
rect 189 194 194 196
rect 196 194 207 196
rect 185 192 207 194
rect 211 196 217 198
rect 211 194 213 196
rect 215 194 217 196
rect 211 192 217 194
rect 130 189 136 191
rect 130 187 132 189
rect 134 187 136 189
rect 130 185 136 187
rect 134 182 136 185
rect 167 183 169 192
rect 178 189 180 192
rect 185 189 187 192
rect 205 189 207 192
rect 215 189 217 192
rect 225 197 227 199
rect 229 197 231 199
rect 225 195 231 197
rect 104 170 106 175
rect 114 170 116 175
rect 66 165 68 169
rect 77 165 79 169
rect 84 165 86 169
rect 124 167 126 172
rect 225 182 227 195
rect 235 191 237 204
rect 307 226 309 231
rect 314 226 316 231
rect 337 229 339 233
rect 369 229 371 233
rect 324 217 326 222
rect 324 201 326 204
rect 269 198 271 201
rect 279 198 281 201
rect 289 198 291 201
rect 307 198 309 201
rect 314 198 316 201
rect 324 199 333 201
rect 267 196 273 198
rect 267 194 269 196
rect 271 194 273 196
rect 267 192 273 194
rect 277 196 283 198
rect 277 194 279 196
rect 281 194 283 196
rect 277 192 283 194
rect 287 196 309 198
rect 287 194 289 196
rect 291 194 296 196
rect 298 194 309 196
rect 287 192 309 194
rect 313 196 319 198
rect 313 194 315 196
rect 317 194 319 196
rect 313 192 319 194
rect 231 189 237 191
rect 231 187 233 189
rect 235 187 237 189
rect 231 185 237 187
rect 235 182 237 185
rect 269 183 271 192
rect 280 189 282 192
rect 287 189 289 192
rect 307 189 309 192
rect 317 189 319 192
rect 327 197 329 199
rect 331 197 333 199
rect 327 195 333 197
rect 205 170 207 175
rect 215 170 217 175
rect 134 165 136 169
rect 167 165 169 169
rect 178 165 180 169
rect 185 165 187 169
rect 225 167 227 172
rect 327 182 329 195
rect 337 191 339 204
rect 382 229 384 233
rect 389 229 391 233
rect 422 229 424 233
rect 432 229 434 233
rect 442 229 444 233
rect 460 226 462 231
rect 467 226 469 231
rect 490 229 492 233
rect 523 229 525 233
rect 533 229 535 233
rect 543 229 545 233
rect 477 217 479 222
rect 477 201 479 204
rect 333 189 339 191
rect 369 198 371 201
rect 382 198 384 201
rect 389 198 391 201
rect 422 198 424 201
rect 432 198 434 201
rect 442 198 444 201
rect 460 198 462 201
rect 467 198 469 201
rect 477 199 486 201
rect 369 196 375 198
rect 369 194 371 196
rect 373 194 375 196
rect 369 192 375 194
rect 379 196 385 198
rect 379 194 381 196
rect 383 194 385 196
rect 379 192 385 194
rect 389 196 398 198
rect 389 194 394 196
rect 396 194 398 196
rect 389 192 398 194
rect 420 196 426 198
rect 420 194 422 196
rect 424 194 426 196
rect 420 192 426 194
rect 430 196 436 198
rect 430 194 432 196
rect 434 194 436 196
rect 430 192 436 194
rect 440 196 462 198
rect 440 194 442 196
rect 444 194 449 196
rect 451 194 462 196
rect 440 192 462 194
rect 466 196 472 198
rect 466 194 468 196
rect 470 194 472 196
rect 466 192 472 194
rect 369 189 371 192
rect 333 187 335 189
rect 337 187 339 189
rect 333 185 339 187
rect 337 182 339 185
rect 307 170 309 175
rect 317 170 319 175
rect 235 165 237 169
rect 269 165 271 169
rect 280 165 282 169
rect 287 165 289 169
rect 327 167 329 172
rect 379 184 381 192
rect 389 186 391 192
rect 422 183 424 192
rect 433 189 435 192
rect 440 189 442 192
rect 460 189 462 192
rect 470 189 472 192
rect 480 197 482 199
rect 484 197 486 199
rect 480 195 486 197
rect 369 170 371 175
rect 379 171 381 176
rect 389 174 391 178
rect 337 165 339 169
rect 480 182 482 195
rect 490 191 492 204
rect 561 226 563 231
rect 568 226 570 231
rect 591 229 593 233
rect 622 229 624 233
rect 632 229 634 233
rect 642 229 644 233
rect 578 217 580 222
rect 578 201 580 204
rect 523 198 525 201
rect 533 198 535 201
rect 543 198 545 201
rect 561 198 563 201
rect 568 198 570 201
rect 578 199 587 201
rect 521 196 527 198
rect 521 194 523 196
rect 525 194 527 196
rect 521 192 527 194
rect 531 196 537 198
rect 531 194 533 196
rect 535 194 537 196
rect 531 192 537 194
rect 541 196 563 198
rect 541 194 543 196
rect 545 194 550 196
rect 552 194 563 196
rect 541 192 563 194
rect 567 196 573 198
rect 567 194 569 196
rect 571 194 573 196
rect 567 192 573 194
rect 486 189 492 191
rect 486 187 488 189
rect 490 187 492 189
rect 486 185 492 187
rect 490 182 492 185
rect 523 183 525 192
rect 534 189 536 192
rect 541 189 543 192
rect 561 189 563 192
rect 571 189 573 192
rect 581 197 583 199
rect 585 197 587 199
rect 581 195 587 197
rect 460 170 462 175
rect 470 170 472 175
rect 422 165 424 169
rect 433 165 435 169
rect 440 165 442 169
rect 480 167 482 172
rect 581 182 583 195
rect 591 191 593 204
rect 660 226 662 231
rect 667 226 669 231
rect 690 229 692 233
rect 677 217 679 222
rect 677 201 679 204
rect 622 198 624 201
rect 632 198 634 201
rect 642 198 644 201
rect 660 198 662 201
rect 667 198 669 201
rect 677 199 686 201
rect 620 196 626 198
rect 620 194 622 196
rect 624 194 626 196
rect 620 192 626 194
rect 630 196 636 198
rect 630 194 632 196
rect 634 194 636 196
rect 630 192 636 194
rect 640 196 662 198
rect 640 194 642 196
rect 644 194 649 196
rect 651 194 662 196
rect 640 192 662 194
rect 666 196 672 198
rect 666 194 668 196
rect 670 194 672 196
rect 666 192 672 194
rect 587 189 593 191
rect 587 187 589 189
rect 591 187 593 189
rect 587 185 593 187
rect 591 182 593 185
rect 622 183 624 192
rect 633 189 635 192
rect 640 189 642 192
rect 660 189 662 192
rect 670 189 672 192
rect 680 197 682 199
rect 684 197 686 199
rect 680 195 686 197
rect 561 170 563 175
rect 571 170 573 175
rect 490 165 492 169
rect 523 165 525 169
rect 534 165 536 169
rect 541 165 543 169
rect 581 167 583 172
rect 680 182 682 195
rect 690 191 692 204
rect 686 189 692 191
rect 686 187 688 189
rect 690 187 692 189
rect 686 185 692 187
rect 690 182 692 185
rect 660 170 662 175
rect 670 170 672 175
rect 591 165 593 169
rect 622 165 624 169
rect 633 165 635 169
rect 640 165 642 169
rect 680 167 682 172
rect 690 165 692 169
rect 27 157 29 161
rect 38 157 40 161
rect 45 157 47 161
rect 27 134 29 143
rect 65 151 67 156
rect 75 151 77 156
rect 85 154 87 159
rect 95 157 97 161
rect 168 157 170 161
rect 179 157 181 161
rect 186 157 188 161
rect 115 151 117 156
rect 38 134 40 137
rect 45 134 47 137
rect 65 134 67 137
rect 75 134 77 137
rect 25 132 31 134
rect 25 130 27 132
rect 29 130 31 132
rect 25 128 31 130
rect 35 132 41 134
rect 35 130 37 132
rect 39 130 41 132
rect 35 128 41 130
rect 45 132 67 134
rect 45 130 47 132
rect 49 130 54 132
rect 56 130 67 132
rect 45 128 67 130
rect 71 132 77 134
rect 71 130 73 132
rect 75 130 77 132
rect 71 128 77 130
rect 85 131 87 144
rect 95 141 97 144
rect 91 139 97 141
rect 91 137 93 139
rect 95 137 97 139
rect 125 150 127 155
rect 135 148 137 152
rect 91 135 97 137
rect 85 129 91 131
rect 27 125 29 128
rect 37 125 39 128
rect 47 125 49 128
rect 65 125 67 128
rect 72 125 74 128
rect 85 127 87 129
rect 89 127 91 129
rect 82 125 91 127
rect 82 122 84 125
rect 95 122 97 135
rect 115 134 117 137
rect 125 134 127 142
rect 135 134 137 140
rect 168 134 170 143
rect 206 151 208 156
rect 216 151 218 156
rect 226 154 228 159
rect 236 157 238 161
rect 268 157 270 161
rect 278 154 280 159
rect 318 157 320 161
rect 325 157 327 161
rect 336 157 338 161
rect 288 151 290 156
rect 298 151 300 156
rect 179 134 181 137
rect 186 134 188 137
rect 206 134 208 137
rect 216 134 218 137
rect 115 132 121 134
rect 115 130 117 132
rect 119 130 121 132
rect 115 128 121 130
rect 125 132 131 134
rect 125 130 127 132
rect 129 130 131 132
rect 125 128 131 130
rect 135 132 144 134
rect 135 130 140 132
rect 142 130 144 132
rect 135 128 144 130
rect 166 132 172 134
rect 166 130 168 132
rect 170 130 172 132
rect 166 128 172 130
rect 176 132 182 134
rect 176 130 178 132
rect 180 130 182 132
rect 176 128 182 130
rect 186 132 208 134
rect 186 130 188 132
rect 190 130 195 132
rect 197 130 208 132
rect 186 128 208 130
rect 212 132 218 134
rect 212 130 214 132
rect 216 130 218 132
rect 212 128 218 130
rect 226 131 228 144
rect 236 141 238 144
rect 232 139 238 141
rect 232 137 234 139
rect 236 137 238 139
rect 232 135 238 137
rect 226 129 232 131
rect 115 125 117 128
rect 128 125 130 128
rect 135 125 137 128
rect 168 125 170 128
rect 178 125 180 128
rect 188 125 190 128
rect 206 125 208 128
rect 213 125 215 128
rect 226 127 228 129
rect 230 127 232 129
rect 223 125 232 127
rect 82 104 84 109
rect 27 93 29 97
rect 37 93 39 97
rect 47 93 49 97
rect 65 95 67 100
rect 72 95 74 100
rect 95 93 97 97
rect 115 93 117 97
rect 223 122 225 125
rect 236 122 238 135
rect 268 141 270 144
rect 268 139 274 141
rect 268 137 270 139
rect 272 137 274 139
rect 268 135 274 137
rect 268 122 270 135
rect 278 131 280 144
rect 422 157 424 161
rect 433 157 435 161
rect 440 157 442 161
rect 369 151 371 156
rect 274 129 280 131
rect 274 127 276 129
rect 278 127 280 129
rect 288 134 290 137
rect 298 134 300 137
rect 318 134 320 137
rect 325 134 327 137
rect 336 134 338 143
rect 379 150 381 155
rect 389 148 391 152
rect 369 134 371 137
rect 379 134 381 142
rect 389 134 391 140
rect 422 134 424 143
rect 460 151 462 156
rect 470 151 472 156
rect 480 154 482 159
rect 490 157 492 161
rect 523 157 525 161
rect 534 157 536 161
rect 541 157 543 161
rect 433 134 435 137
rect 440 134 442 137
rect 460 134 462 137
rect 470 134 472 137
rect 288 132 294 134
rect 288 130 290 132
rect 292 130 294 132
rect 288 128 294 130
rect 298 132 320 134
rect 298 130 309 132
rect 311 130 316 132
rect 318 130 320 132
rect 298 128 320 130
rect 324 132 330 134
rect 324 130 326 132
rect 328 130 330 132
rect 324 128 330 130
rect 334 132 340 134
rect 334 130 336 132
rect 338 130 340 132
rect 334 128 340 130
rect 369 132 375 134
rect 369 130 371 132
rect 373 130 375 132
rect 369 128 375 130
rect 379 132 385 134
rect 379 130 381 132
rect 383 130 385 132
rect 379 128 385 130
rect 389 132 398 134
rect 389 130 394 132
rect 396 130 398 132
rect 389 128 398 130
rect 420 132 426 134
rect 420 130 422 132
rect 424 130 426 132
rect 420 128 426 130
rect 430 132 436 134
rect 430 130 432 132
rect 434 130 436 132
rect 430 128 436 130
rect 440 132 462 134
rect 440 130 442 132
rect 444 130 449 132
rect 451 130 462 132
rect 440 128 462 130
rect 466 132 472 134
rect 466 130 468 132
rect 470 130 472 132
rect 466 128 472 130
rect 480 131 482 144
rect 490 141 492 144
rect 486 139 492 141
rect 486 137 488 139
rect 490 137 492 139
rect 486 135 492 137
rect 480 129 486 131
rect 274 125 283 127
rect 291 125 293 128
rect 298 125 300 128
rect 316 125 318 128
rect 326 125 328 128
rect 336 125 338 128
rect 369 125 371 128
rect 382 125 384 128
rect 389 125 391 128
rect 422 125 424 128
rect 432 125 434 128
rect 442 125 444 128
rect 460 125 462 128
rect 467 125 469 128
rect 480 127 482 129
rect 484 127 486 129
rect 477 125 486 127
rect 281 122 283 125
rect 223 104 225 109
rect 128 93 130 97
rect 135 93 137 97
rect 168 93 170 97
rect 178 93 180 97
rect 188 93 190 97
rect 206 95 208 100
rect 213 95 215 100
rect 281 104 283 109
rect 236 93 238 97
rect 268 93 270 97
rect 291 95 293 100
rect 298 95 300 100
rect 316 93 318 97
rect 326 93 328 97
rect 336 93 338 97
rect 369 93 371 97
rect 477 122 479 125
rect 490 122 492 135
rect 523 134 525 143
rect 561 151 563 156
rect 571 151 573 156
rect 581 154 583 159
rect 591 157 593 161
rect 622 157 624 161
rect 633 157 635 161
rect 640 157 642 161
rect 534 134 536 137
rect 541 134 543 137
rect 561 134 563 137
rect 571 134 573 137
rect 521 132 527 134
rect 521 130 523 132
rect 525 130 527 132
rect 521 128 527 130
rect 531 132 537 134
rect 531 130 533 132
rect 535 130 537 132
rect 531 128 537 130
rect 541 132 563 134
rect 541 130 543 132
rect 545 130 550 132
rect 552 130 563 132
rect 541 128 563 130
rect 567 132 573 134
rect 567 130 569 132
rect 571 130 573 132
rect 567 128 573 130
rect 581 131 583 144
rect 591 141 593 144
rect 587 139 593 141
rect 587 137 589 139
rect 591 137 593 139
rect 587 135 593 137
rect 581 129 587 131
rect 523 125 525 128
rect 533 125 535 128
rect 543 125 545 128
rect 561 125 563 128
rect 568 125 570 128
rect 581 127 583 129
rect 585 127 587 129
rect 578 125 587 127
rect 477 104 479 109
rect 382 93 384 97
rect 389 93 391 97
rect 422 93 424 97
rect 432 93 434 97
rect 442 93 444 97
rect 460 95 462 100
rect 467 95 469 100
rect 578 122 580 125
rect 591 122 593 135
rect 622 134 624 143
rect 660 151 662 156
rect 670 151 672 156
rect 680 154 682 159
rect 690 157 692 161
rect 633 134 635 137
rect 640 134 642 137
rect 660 134 662 137
rect 670 134 672 137
rect 620 132 626 134
rect 620 130 622 132
rect 624 130 626 132
rect 620 128 626 130
rect 630 132 636 134
rect 630 130 632 132
rect 634 130 636 132
rect 630 128 636 130
rect 640 132 662 134
rect 640 130 642 132
rect 644 130 649 132
rect 651 130 662 132
rect 640 128 662 130
rect 666 132 672 134
rect 666 130 668 132
rect 670 130 672 132
rect 666 128 672 130
rect 680 131 682 144
rect 690 141 692 144
rect 686 139 692 141
rect 686 137 688 139
rect 690 137 692 139
rect 686 135 692 137
rect 680 129 686 131
rect 622 125 624 128
rect 632 125 634 128
rect 642 125 644 128
rect 660 125 662 128
rect 667 125 669 128
rect 680 127 682 129
rect 684 127 686 129
rect 677 125 686 127
rect 578 104 580 109
rect 490 93 492 97
rect 523 93 525 97
rect 533 93 535 97
rect 543 93 545 97
rect 561 95 563 100
rect 568 95 570 100
rect 677 122 679 125
rect 690 122 692 135
rect 677 104 679 109
rect 591 93 593 97
rect 622 93 624 97
rect 632 93 634 97
rect 642 93 644 97
rect 660 95 662 100
rect 667 95 669 100
rect 690 93 692 97
rect 25 85 27 89
rect 38 85 40 89
rect 45 85 47 89
rect 66 85 68 89
rect 76 85 78 89
rect 86 85 88 89
rect 104 82 106 87
rect 111 82 113 87
rect 134 85 136 89
rect 167 85 169 89
rect 177 85 179 89
rect 187 85 189 89
rect 121 73 123 78
rect 121 57 123 60
rect 25 54 27 57
rect 38 54 40 57
rect 45 54 47 57
rect 66 54 68 57
rect 76 54 78 57
rect 86 54 88 57
rect 104 54 106 57
rect 111 54 113 57
rect 121 55 130 57
rect 25 52 31 54
rect 25 50 27 52
rect 29 50 31 52
rect 25 48 31 50
rect 35 52 41 54
rect 35 50 37 52
rect 39 50 41 52
rect 35 48 41 50
rect 45 52 54 54
rect 45 50 50 52
rect 52 50 54 52
rect 45 48 54 50
rect 64 52 70 54
rect 64 50 66 52
rect 68 50 70 52
rect 64 48 70 50
rect 74 52 80 54
rect 74 50 76 52
rect 78 50 80 52
rect 74 48 80 50
rect 84 52 106 54
rect 84 50 86 52
rect 88 50 93 52
rect 95 50 106 52
rect 84 48 106 50
rect 110 52 116 54
rect 110 50 112 52
rect 114 50 116 52
rect 110 48 116 50
rect 25 45 27 48
rect 35 40 37 48
rect 45 42 47 48
rect 66 39 68 48
rect 77 45 79 48
rect 84 45 86 48
rect 104 45 106 48
rect 114 45 116 48
rect 124 53 126 55
rect 128 53 130 55
rect 124 51 130 53
rect 25 26 27 31
rect 35 27 37 32
rect 45 30 47 34
rect 124 38 126 51
rect 134 47 136 60
rect 205 82 207 87
rect 212 82 214 87
rect 235 85 237 89
rect 268 85 270 89
rect 278 85 280 89
rect 288 85 290 89
rect 222 73 224 78
rect 222 57 224 60
rect 167 54 169 57
rect 177 54 179 57
rect 187 54 189 57
rect 205 54 207 57
rect 212 54 214 57
rect 222 55 231 57
rect 165 52 171 54
rect 165 50 167 52
rect 169 50 171 52
rect 165 48 171 50
rect 175 52 181 54
rect 175 50 177 52
rect 179 50 181 52
rect 175 48 181 50
rect 185 52 207 54
rect 185 50 187 52
rect 189 50 194 52
rect 196 50 207 52
rect 185 48 207 50
rect 211 52 217 54
rect 211 50 213 52
rect 215 50 217 52
rect 211 48 217 50
rect 130 45 136 47
rect 130 43 132 45
rect 134 43 136 45
rect 130 41 136 43
rect 134 38 136 41
rect 167 39 169 48
rect 178 45 180 48
rect 185 45 187 48
rect 205 45 207 48
rect 215 45 217 48
rect 225 53 227 55
rect 229 53 231 55
rect 225 51 231 53
rect 104 26 106 31
rect 114 26 116 31
rect 66 21 68 25
rect 77 21 79 25
rect 84 21 86 25
rect 124 23 126 28
rect 225 38 227 51
rect 235 47 237 60
rect 306 82 308 87
rect 313 82 315 87
rect 336 85 338 89
rect 368 85 370 89
rect 323 73 325 78
rect 323 57 325 60
rect 268 54 270 57
rect 278 54 280 57
rect 288 54 290 57
rect 306 54 308 57
rect 313 54 315 57
rect 323 55 332 57
rect 266 52 272 54
rect 266 50 268 52
rect 270 50 272 52
rect 266 48 272 50
rect 276 52 282 54
rect 276 50 278 52
rect 280 50 282 52
rect 276 48 282 50
rect 286 52 308 54
rect 286 50 288 52
rect 290 50 295 52
rect 297 50 308 52
rect 286 48 308 50
rect 312 52 318 54
rect 312 50 314 52
rect 316 50 318 52
rect 312 48 318 50
rect 231 45 237 47
rect 231 43 233 45
rect 235 43 237 45
rect 231 41 237 43
rect 235 38 237 41
rect 268 39 270 48
rect 279 45 281 48
rect 286 45 288 48
rect 306 45 308 48
rect 316 45 318 48
rect 326 53 328 55
rect 330 53 332 55
rect 326 51 332 53
rect 205 26 207 31
rect 215 26 217 31
rect 134 21 136 25
rect 167 21 169 25
rect 178 21 180 25
rect 185 21 187 25
rect 225 23 227 28
rect 326 38 328 51
rect 336 47 338 60
rect 381 85 383 89
rect 388 85 390 89
rect 421 85 423 89
rect 431 85 433 89
rect 441 85 443 89
rect 459 82 461 87
rect 466 82 468 87
rect 489 85 491 89
rect 522 85 524 89
rect 532 85 534 89
rect 542 85 544 89
rect 476 73 478 78
rect 476 57 478 60
rect 332 45 338 47
rect 368 54 370 57
rect 381 54 383 57
rect 388 54 390 57
rect 421 54 423 57
rect 431 54 433 57
rect 441 54 443 57
rect 459 54 461 57
rect 466 54 468 57
rect 476 55 485 57
rect 368 52 374 54
rect 368 50 370 52
rect 372 50 374 52
rect 368 48 374 50
rect 378 52 384 54
rect 378 50 380 52
rect 382 50 384 52
rect 378 48 384 50
rect 388 52 397 54
rect 388 50 393 52
rect 395 50 397 52
rect 388 48 397 50
rect 419 52 425 54
rect 419 50 421 52
rect 423 50 425 52
rect 419 48 425 50
rect 429 52 435 54
rect 429 50 431 52
rect 433 50 435 52
rect 429 48 435 50
rect 439 52 461 54
rect 439 50 441 52
rect 443 50 448 52
rect 450 50 461 52
rect 439 48 461 50
rect 465 52 471 54
rect 465 50 467 52
rect 469 50 471 52
rect 465 48 471 50
rect 368 45 370 48
rect 332 43 334 45
rect 336 43 338 45
rect 332 41 338 43
rect 336 38 338 41
rect 306 26 308 31
rect 316 26 318 31
rect 235 21 237 25
rect 268 21 270 25
rect 279 21 281 25
rect 286 21 288 25
rect 326 23 328 28
rect 378 40 380 48
rect 388 42 390 48
rect 421 39 423 48
rect 432 45 434 48
rect 439 45 441 48
rect 459 45 461 48
rect 469 45 471 48
rect 479 53 481 55
rect 483 53 485 55
rect 479 51 485 53
rect 368 26 370 31
rect 378 27 380 32
rect 388 30 390 34
rect 336 21 338 25
rect 479 38 481 51
rect 489 47 491 60
rect 560 82 562 87
rect 567 82 569 87
rect 590 85 592 89
rect 621 85 623 89
rect 631 85 633 89
rect 641 85 643 89
rect 577 73 579 78
rect 577 57 579 60
rect 522 54 524 57
rect 532 54 534 57
rect 542 54 544 57
rect 560 54 562 57
rect 567 54 569 57
rect 577 55 586 57
rect 520 52 526 54
rect 520 50 522 52
rect 524 50 526 52
rect 520 48 526 50
rect 530 52 536 54
rect 530 50 532 52
rect 534 50 536 52
rect 530 48 536 50
rect 540 52 562 54
rect 540 50 542 52
rect 544 50 549 52
rect 551 50 562 52
rect 540 48 562 50
rect 566 52 572 54
rect 566 50 568 52
rect 570 50 572 52
rect 566 48 572 50
rect 485 45 491 47
rect 485 43 487 45
rect 489 43 491 45
rect 485 41 491 43
rect 489 38 491 41
rect 522 39 524 48
rect 533 45 535 48
rect 540 45 542 48
rect 560 45 562 48
rect 570 45 572 48
rect 580 53 582 55
rect 584 53 586 55
rect 580 51 586 53
rect 459 26 461 31
rect 469 26 471 31
rect 421 21 423 25
rect 432 21 434 25
rect 439 21 441 25
rect 479 23 481 28
rect 580 38 582 51
rect 590 47 592 60
rect 659 82 661 87
rect 666 82 668 87
rect 689 85 691 89
rect 676 73 678 78
rect 676 57 678 60
rect 621 54 623 57
rect 631 54 633 57
rect 641 54 643 57
rect 659 54 661 57
rect 666 54 668 57
rect 676 55 685 57
rect 619 52 625 54
rect 619 50 621 52
rect 623 50 625 52
rect 619 48 625 50
rect 629 52 635 54
rect 629 50 631 52
rect 633 50 635 52
rect 629 48 635 50
rect 639 52 661 54
rect 639 50 641 52
rect 643 50 648 52
rect 650 50 661 52
rect 639 48 661 50
rect 665 52 671 54
rect 665 50 667 52
rect 669 50 671 52
rect 665 48 671 50
rect 586 45 592 47
rect 586 43 588 45
rect 590 43 592 45
rect 586 41 592 43
rect 590 38 592 41
rect 621 39 623 48
rect 632 45 634 48
rect 639 45 641 48
rect 659 45 661 48
rect 669 45 671 48
rect 679 53 681 55
rect 683 53 685 55
rect 679 51 685 53
rect 560 26 562 31
rect 570 26 572 31
rect 489 21 491 25
rect 522 21 524 25
rect 533 21 535 25
rect 540 21 542 25
rect 580 23 582 28
rect 679 38 681 51
rect 689 47 691 60
rect 685 45 691 47
rect 685 43 687 45
rect 689 43 691 45
rect 685 41 691 43
rect 689 38 691 41
rect 659 26 661 31
rect 669 26 671 31
rect 590 21 592 25
rect 621 21 623 25
rect 632 21 634 25
rect 639 21 641 25
rect 679 23 681 28
rect 689 21 691 25
<< ndif >>
rect 20 326 25 333
rect 18 324 25 326
rect 18 322 20 324
rect 22 322 25 324
rect 18 320 25 322
rect 27 320 32 333
rect 34 320 45 333
rect 36 319 45 320
rect 47 331 54 333
rect 47 329 50 331
rect 52 329 54 331
rect 47 323 54 329
rect 60 326 65 333
rect 47 321 50 323
rect 52 321 54 323
rect 47 319 54 321
rect 58 324 65 326
rect 58 322 60 324
rect 62 322 65 324
rect 58 320 65 322
rect 67 320 72 333
rect 74 320 85 333
rect 36 314 43 319
rect 76 319 85 320
rect 87 331 94 333
rect 87 329 90 331
rect 92 329 94 331
rect 87 323 94 329
rect 110 327 117 333
rect 87 321 90 323
rect 92 321 94 323
rect 87 319 94 321
rect 99 324 106 327
rect 99 322 101 324
rect 103 322 106 324
rect 99 320 106 322
rect 76 314 83 319
rect 36 312 39 314
rect 41 312 43 314
rect 36 310 43 312
rect 76 312 79 314
rect 81 312 83 314
rect 101 313 106 320
rect 108 317 117 327
rect 108 315 112 317
rect 114 315 117 317
rect 108 313 117 315
rect 119 313 124 333
rect 126 326 131 333
rect 137 331 144 333
rect 137 329 139 331
rect 141 329 144 331
rect 126 324 133 326
rect 126 322 129 324
rect 131 322 133 324
rect 126 320 133 322
rect 137 324 144 329
rect 137 322 139 324
rect 141 322 144 324
rect 126 313 131 320
rect 137 319 144 322
rect 146 331 154 333
rect 146 329 149 331
rect 151 329 154 331
rect 146 319 154 329
rect 156 326 161 333
rect 217 326 222 333
rect 156 323 164 326
rect 156 321 159 323
rect 161 321 164 323
rect 156 319 164 321
rect 159 316 164 319
rect 166 320 174 326
rect 166 318 169 320
rect 171 318 174 320
rect 166 316 174 318
rect 76 310 83 312
rect 169 313 174 316
rect 176 324 183 326
rect 176 322 179 324
rect 181 322 183 324
rect 176 320 183 322
rect 195 324 202 326
rect 195 322 197 324
rect 199 322 202 324
rect 195 320 202 322
rect 176 313 181 320
rect 197 313 202 320
rect 204 320 212 326
rect 204 318 207 320
rect 209 318 212 320
rect 204 316 212 318
rect 214 323 222 326
rect 214 321 217 323
rect 219 321 222 323
rect 214 319 222 321
rect 224 331 232 333
rect 224 329 227 331
rect 229 329 232 331
rect 224 319 232 329
rect 234 331 241 333
rect 234 329 237 331
rect 239 329 241 331
rect 234 324 241 329
rect 247 326 252 333
rect 234 322 237 324
rect 239 322 241 324
rect 234 319 241 322
rect 245 324 252 326
rect 245 322 247 324
rect 249 322 252 324
rect 245 320 252 322
rect 214 316 219 319
rect 204 313 209 316
rect 247 313 252 320
rect 254 313 259 333
rect 261 327 268 333
rect 284 331 291 333
rect 284 329 286 331
rect 288 329 291 331
rect 261 317 270 327
rect 261 315 264 317
rect 266 315 270 317
rect 261 313 270 315
rect 272 324 279 327
rect 272 322 275 324
rect 277 322 279 324
rect 272 320 279 322
rect 284 323 291 329
rect 284 321 286 323
rect 288 321 291 323
rect 272 313 277 320
rect 284 319 291 321
rect 293 320 304 333
rect 306 320 311 333
rect 313 326 318 333
rect 324 331 331 333
rect 324 329 326 331
rect 328 329 331 331
rect 313 324 320 326
rect 313 322 316 324
rect 318 322 320 324
rect 313 320 320 322
rect 324 323 331 329
rect 324 321 326 323
rect 328 321 331 323
rect 293 319 302 320
rect 295 314 302 319
rect 324 319 331 321
rect 333 320 344 333
rect 346 320 351 333
rect 353 326 358 333
rect 387 326 392 333
rect 353 324 360 326
rect 353 322 356 324
rect 358 322 360 324
rect 353 320 360 322
rect 365 324 372 326
rect 365 322 367 324
rect 369 322 372 324
rect 365 320 372 322
rect 333 319 342 320
rect 335 314 342 319
rect 295 312 297 314
rect 299 312 302 314
rect 295 310 302 312
rect 335 312 337 314
rect 339 312 342 314
rect 367 313 372 320
rect 374 320 382 326
rect 374 318 377 320
rect 379 318 382 320
rect 374 316 382 318
rect 384 323 392 326
rect 384 321 387 323
rect 389 321 392 323
rect 384 319 392 321
rect 394 331 402 333
rect 394 329 397 331
rect 399 329 402 331
rect 394 319 402 329
rect 404 331 411 333
rect 404 329 407 331
rect 409 329 411 331
rect 404 324 411 329
rect 417 326 422 333
rect 404 322 407 324
rect 409 322 411 324
rect 404 319 411 322
rect 415 324 422 326
rect 415 322 417 324
rect 419 322 422 324
rect 415 320 422 322
rect 384 316 389 319
rect 374 313 379 316
rect 335 310 342 312
rect 417 313 422 320
rect 424 313 429 333
rect 431 327 438 333
rect 454 331 461 333
rect 454 329 456 331
rect 458 329 461 331
rect 431 317 440 327
rect 431 315 434 317
rect 436 315 440 317
rect 431 313 440 315
rect 442 324 449 327
rect 442 322 445 324
rect 447 322 449 324
rect 442 320 449 322
rect 454 323 461 329
rect 454 321 456 323
rect 458 321 461 323
rect 442 313 447 320
rect 454 319 461 321
rect 463 320 474 333
rect 476 320 481 333
rect 483 326 488 333
rect 494 331 501 333
rect 494 329 496 331
rect 498 329 501 331
rect 483 324 490 326
rect 483 322 486 324
rect 488 322 490 324
rect 483 320 490 322
rect 494 323 501 329
rect 494 321 496 323
rect 498 321 501 323
rect 463 319 472 320
rect 465 314 472 319
rect 494 319 501 321
rect 503 320 514 333
rect 516 320 521 333
rect 523 326 528 333
rect 536 326 541 333
rect 523 324 530 326
rect 523 322 526 324
rect 528 322 530 324
rect 523 320 530 322
rect 534 324 541 326
rect 534 322 536 324
rect 538 322 541 324
rect 534 320 541 322
rect 543 320 548 333
rect 550 320 561 333
rect 503 319 512 320
rect 505 314 512 319
rect 552 319 561 320
rect 563 331 570 333
rect 563 329 566 331
rect 568 329 570 331
rect 563 323 570 329
rect 576 326 581 333
rect 563 321 566 323
rect 568 321 570 323
rect 563 319 570 321
rect 574 324 581 326
rect 574 322 576 324
rect 578 322 581 324
rect 574 320 581 322
rect 583 320 588 333
rect 590 320 601 333
rect 465 312 467 314
rect 469 312 472 314
rect 465 310 472 312
rect 505 312 507 314
rect 509 312 512 314
rect 505 310 512 312
rect 552 314 559 319
rect 592 319 601 320
rect 603 331 610 333
rect 603 329 606 331
rect 608 329 610 331
rect 603 323 610 329
rect 626 327 633 333
rect 603 321 606 323
rect 608 321 610 323
rect 603 319 610 321
rect 615 324 622 327
rect 615 322 617 324
rect 619 322 622 324
rect 615 320 622 322
rect 592 314 599 319
rect 552 312 555 314
rect 557 312 559 314
rect 552 310 559 312
rect 592 312 595 314
rect 597 312 599 314
rect 617 313 622 320
rect 624 317 633 327
rect 624 315 628 317
rect 630 315 633 317
rect 624 313 633 315
rect 635 313 640 333
rect 642 326 647 333
rect 653 331 660 333
rect 653 329 655 331
rect 657 329 660 331
rect 642 324 649 326
rect 642 322 645 324
rect 647 322 649 324
rect 642 320 649 322
rect 653 324 660 329
rect 653 322 655 324
rect 657 322 660 324
rect 642 313 647 320
rect 653 319 660 322
rect 662 331 670 333
rect 662 329 665 331
rect 667 329 670 331
rect 662 319 670 329
rect 672 326 677 333
rect 672 323 680 326
rect 672 321 675 323
rect 677 321 680 323
rect 672 319 680 321
rect 675 316 680 319
rect 682 320 690 326
rect 682 318 685 320
rect 687 318 690 320
rect 682 316 690 318
rect 592 310 599 312
rect 685 313 690 316
rect 692 324 699 326
rect 692 322 695 324
rect 697 322 699 324
rect 692 320 699 322
rect 692 313 697 320
rect 36 302 43 304
rect 36 300 39 302
rect 41 300 43 302
rect 76 302 83 304
rect 76 300 79 302
rect 81 300 83 302
rect 36 295 43 300
rect 36 294 45 295
rect 18 292 25 294
rect 18 290 20 292
rect 22 290 25 292
rect 18 288 25 290
rect 20 281 25 288
rect 27 281 32 294
rect 34 281 45 294
rect 47 293 54 295
rect 76 295 83 300
rect 76 294 85 295
rect 47 291 50 293
rect 52 291 54 293
rect 47 285 54 291
rect 58 292 65 294
rect 58 290 60 292
rect 62 290 65 292
rect 58 288 65 290
rect 47 283 50 285
rect 52 283 54 285
rect 47 281 54 283
rect 60 281 65 288
rect 67 281 72 294
rect 74 281 85 294
rect 87 293 94 295
rect 101 294 106 301
rect 87 291 90 293
rect 92 291 94 293
rect 87 285 94 291
rect 99 292 106 294
rect 99 290 101 292
rect 103 290 106 292
rect 99 287 106 290
rect 108 299 117 301
rect 108 297 112 299
rect 114 297 117 299
rect 108 287 117 297
rect 87 283 90 285
rect 92 283 94 285
rect 87 281 94 283
rect 110 281 117 287
rect 119 281 124 301
rect 126 294 131 301
rect 169 298 174 301
rect 159 295 164 298
rect 126 292 133 294
rect 126 290 129 292
rect 131 290 133 292
rect 126 288 133 290
rect 137 292 144 295
rect 137 290 139 292
rect 141 290 144 292
rect 126 281 131 288
rect 137 285 144 290
rect 137 283 139 285
rect 141 283 144 285
rect 137 281 144 283
rect 146 285 154 295
rect 146 283 149 285
rect 151 283 154 285
rect 146 281 154 283
rect 156 293 164 295
rect 156 291 159 293
rect 161 291 164 293
rect 156 288 164 291
rect 166 296 174 298
rect 166 294 169 296
rect 171 294 174 296
rect 166 288 174 294
rect 176 294 181 301
rect 197 294 202 301
rect 176 292 183 294
rect 176 290 179 292
rect 181 290 183 292
rect 176 288 183 290
rect 195 292 202 294
rect 195 290 197 292
rect 199 290 202 292
rect 195 288 202 290
rect 204 298 209 301
rect 295 302 302 304
rect 204 296 212 298
rect 204 294 207 296
rect 209 294 212 296
rect 204 288 212 294
rect 214 295 219 298
rect 214 293 222 295
rect 214 291 217 293
rect 219 291 222 293
rect 214 288 222 291
rect 156 281 161 288
rect 217 281 222 288
rect 224 285 232 295
rect 224 283 227 285
rect 229 283 232 285
rect 224 281 232 283
rect 234 292 241 295
rect 247 294 252 301
rect 234 290 237 292
rect 239 290 241 292
rect 234 285 241 290
rect 245 292 252 294
rect 245 290 247 292
rect 249 290 252 292
rect 245 288 252 290
rect 234 283 237 285
rect 239 283 241 285
rect 234 281 241 283
rect 247 281 252 288
rect 254 281 259 301
rect 261 299 270 301
rect 261 297 264 299
rect 266 297 270 299
rect 261 287 270 297
rect 272 294 277 301
rect 295 300 297 302
rect 299 300 302 302
rect 335 302 342 304
rect 335 300 337 302
rect 339 300 342 302
rect 295 295 302 300
rect 272 292 279 294
rect 272 290 275 292
rect 277 290 279 292
rect 272 287 279 290
rect 284 293 291 295
rect 284 291 286 293
rect 288 291 291 293
rect 261 281 268 287
rect 284 285 291 291
rect 284 283 286 285
rect 288 283 291 285
rect 284 281 291 283
rect 293 294 302 295
rect 335 295 342 300
rect 293 281 304 294
rect 306 281 311 294
rect 313 292 320 294
rect 313 290 316 292
rect 318 290 320 292
rect 313 288 320 290
rect 324 293 331 295
rect 324 291 326 293
rect 328 291 331 293
rect 313 281 318 288
rect 324 285 331 291
rect 324 283 326 285
rect 328 283 331 285
rect 324 281 331 283
rect 333 294 342 295
rect 367 294 372 301
rect 333 281 344 294
rect 346 281 351 294
rect 353 292 360 294
rect 353 290 356 292
rect 358 290 360 292
rect 353 288 360 290
rect 365 292 372 294
rect 365 290 367 292
rect 369 290 372 292
rect 365 288 372 290
rect 374 298 379 301
rect 465 302 472 304
rect 374 296 382 298
rect 374 294 377 296
rect 379 294 382 296
rect 374 288 382 294
rect 384 295 389 298
rect 384 293 392 295
rect 384 291 387 293
rect 389 291 392 293
rect 384 288 392 291
rect 353 281 358 288
rect 387 281 392 288
rect 394 285 402 295
rect 394 283 397 285
rect 399 283 402 285
rect 394 281 402 283
rect 404 292 411 295
rect 417 294 422 301
rect 404 290 407 292
rect 409 290 411 292
rect 404 285 411 290
rect 415 292 422 294
rect 415 290 417 292
rect 419 290 422 292
rect 415 288 422 290
rect 404 283 407 285
rect 409 283 411 285
rect 404 281 411 283
rect 417 281 422 288
rect 424 281 429 301
rect 431 299 440 301
rect 431 297 434 299
rect 436 297 440 299
rect 431 287 440 297
rect 442 294 447 301
rect 465 300 467 302
rect 469 300 472 302
rect 505 302 512 304
rect 505 300 507 302
rect 509 300 512 302
rect 465 295 472 300
rect 442 292 449 294
rect 442 290 445 292
rect 447 290 449 292
rect 442 287 449 290
rect 454 293 461 295
rect 454 291 456 293
rect 458 291 461 293
rect 431 281 438 287
rect 454 285 461 291
rect 454 283 456 285
rect 458 283 461 285
rect 454 281 461 283
rect 463 294 472 295
rect 505 295 512 300
rect 552 302 559 304
rect 552 300 555 302
rect 557 300 559 302
rect 592 302 599 304
rect 592 300 595 302
rect 597 300 599 302
rect 463 281 474 294
rect 476 281 481 294
rect 483 292 490 294
rect 483 290 486 292
rect 488 290 490 292
rect 483 288 490 290
rect 494 293 501 295
rect 494 291 496 293
rect 498 291 501 293
rect 483 281 488 288
rect 494 285 501 291
rect 494 283 496 285
rect 498 283 501 285
rect 494 281 501 283
rect 503 294 512 295
rect 552 295 559 300
rect 552 294 561 295
rect 503 281 514 294
rect 516 281 521 294
rect 523 292 530 294
rect 523 290 526 292
rect 528 290 530 292
rect 523 288 530 290
rect 534 292 541 294
rect 534 290 536 292
rect 538 290 541 292
rect 534 288 541 290
rect 523 281 528 288
rect 536 281 541 288
rect 543 281 548 294
rect 550 281 561 294
rect 563 293 570 295
rect 592 295 599 300
rect 592 294 601 295
rect 563 291 566 293
rect 568 291 570 293
rect 563 285 570 291
rect 574 292 581 294
rect 574 290 576 292
rect 578 290 581 292
rect 574 288 581 290
rect 563 283 566 285
rect 568 283 570 285
rect 563 281 570 283
rect 576 281 581 288
rect 583 281 588 294
rect 590 281 601 294
rect 603 293 610 295
rect 617 294 622 301
rect 603 291 606 293
rect 608 291 610 293
rect 603 285 610 291
rect 615 292 622 294
rect 615 290 617 292
rect 619 290 622 292
rect 615 287 622 290
rect 624 299 633 301
rect 624 297 628 299
rect 630 297 633 299
rect 624 287 633 297
rect 603 283 606 285
rect 608 283 610 285
rect 603 281 610 283
rect 626 281 633 287
rect 635 281 640 301
rect 642 294 647 301
rect 685 298 690 301
rect 675 295 680 298
rect 642 292 649 294
rect 642 290 645 292
rect 647 290 649 292
rect 642 288 649 290
rect 653 292 660 295
rect 653 290 655 292
rect 657 290 660 292
rect 642 281 647 288
rect 653 285 660 290
rect 653 283 655 285
rect 657 283 660 285
rect 653 281 660 283
rect 662 285 670 295
rect 662 283 665 285
rect 667 283 670 285
rect 662 281 670 283
rect 672 293 680 295
rect 672 291 675 293
rect 677 291 680 293
rect 672 288 680 291
rect 682 296 690 298
rect 682 294 685 296
rect 687 294 690 296
rect 682 288 690 294
rect 692 294 697 301
rect 692 292 699 294
rect 692 290 695 292
rect 697 290 699 292
rect 692 288 699 290
rect 672 281 677 288
rect 18 187 25 189
rect 18 185 20 187
rect 22 185 25 187
rect 18 180 25 185
rect 18 178 20 180
rect 22 178 25 180
rect 18 175 25 178
rect 27 184 32 189
rect 40 184 45 186
rect 27 180 35 184
rect 27 178 30 180
rect 32 178 35 180
rect 27 176 35 178
rect 37 182 45 184
rect 37 180 40 182
rect 42 180 45 182
rect 37 178 45 180
rect 47 182 54 186
rect 70 183 77 189
rect 47 180 50 182
rect 52 180 54 182
rect 47 178 54 180
rect 59 180 66 183
rect 59 178 61 180
rect 63 178 66 180
rect 37 176 42 178
rect 27 175 32 176
rect 59 176 66 178
rect 61 169 66 176
rect 68 173 77 183
rect 68 171 72 173
rect 74 171 77 173
rect 68 169 77 171
rect 79 169 84 189
rect 86 182 91 189
rect 97 187 104 189
rect 97 185 99 187
rect 101 185 104 187
rect 86 180 93 182
rect 86 178 89 180
rect 91 178 93 180
rect 86 176 93 178
rect 97 180 104 185
rect 97 178 99 180
rect 101 178 104 180
rect 86 169 91 176
rect 97 175 104 178
rect 106 187 114 189
rect 106 185 109 187
rect 111 185 114 187
rect 106 175 114 185
rect 116 182 121 189
rect 171 183 178 189
rect 116 179 124 182
rect 116 177 119 179
rect 121 177 124 179
rect 116 175 124 177
rect 119 172 124 175
rect 126 176 134 182
rect 126 174 129 176
rect 131 174 134 176
rect 126 172 134 174
rect 129 169 134 172
rect 136 180 143 182
rect 136 178 139 180
rect 141 178 143 180
rect 136 176 143 178
rect 160 180 167 183
rect 160 178 162 180
rect 164 178 167 180
rect 160 176 167 178
rect 136 169 141 176
rect 162 169 167 176
rect 169 173 178 183
rect 169 171 173 173
rect 175 171 178 173
rect 169 169 178 171
rect 180 169 185 189
rect 187 182 192 189
rect 198 187 205 189
rect 198 185 200 187
rect 202 185 205 187
rect 187 180 194 182
rect 187 178 190 180
rect 192 178 194 180
rect 187 176 194 178
rect 198 180 205 185
rect 198 178 200 180
rect 202 178 205 180
rect 187 169 192 176
rect 198 175 205 178
rect 207 187 215 189
rect 207 185 210 187
rect 212 185 215 187
rect 207 175 215 185
rect 217 182 222 189
rect 273 183 280 189
rect 217 179 225 182
rect 217 177 220 179
rect 222 177 225 179
rect 217 175 225 177
rect 220 172 225 175
rect 227 176 235 182
rect 227 174 230 176
rect 232 174 235 176
rect 227 172 235 174
rect 230 169 235 172
rect 237 180 244 182
rect 237 178 240 180
rect 242 178 244 180
rect 237 176 244 178
rect 262 180 269 183
rect 262 178 264 180
rect 266 178 269 180
rect 262 176 269 178
rect 237 169 242 176
rect 264 169 269 176
rect 271 173 280 183
rect 271 171 275 173
rect 277 171 280 173
rect 271 169 280 171
rect 282 169 287 189
rect 289 182 294 189
rect 300 187 307 189
rect 300 185 302 187
rect 304 185 307 187
rect 289 180 296 182
rect 289 178 292 180
rect 294 178 296 180
rect 289 176 296 178
rect 300 180 307 185
rect 300 178 302 180
rect 304 178 307 180
rect 289 169 294 176
rect 300 175 307 178
rect 309 187 317 189
rect 309 185 312 187
rect 314 185 317 187
rect 309 175 317 185
rect 319 182 324 189
rect 362 187 369 189
rect 362 185 364 187
rect 366 185 369 187
rect 319 179 327 182
rect 319 177 322 179
rect 324 177 327 179
rect 319 175 327 177
rect 322 172 327 175
rect 329 176 337 182
rect 329 174 332 176
rect 334 174 337 176
rect 329 172 337 174
rect 332 169 337 172
rect 339 180 346 182
rect 339 178 342 180
rect 344 178 346 180
rect 339 176 346 178
rect 362 180 369 185
rect 362 178 364 180
rect 366 178 369 180
rect 339 169 344 176
rect 362 175 369 178
rect 371 184 376 189
rect 384 184 389 186
rect 371 180 379 184
rect 371 178 374 180
rect 376 178 379 180
rect 371 176 379 178
rect 381 182 389 184
rect 381 180 384 182
rect 386 180 389 182
rect 381 178 389 180
rect 391 182 398 186
rect 426 183 433 189
rect 391 180 394 182
rect 396 180 398 182
rect 391 178 398 180
rect 415 180 422 183
rect 415 178 417 180
rect 419 178 422 180
rect 381 176 386 178
rect 371 175 376 176
rect 415 176 422 178
rect 417 169 422 176
rect 424 173 433 183
rect 424 171 428 173
rect 430 171 433 173
rect 424 169 433 171
rect 435 169 440 189
rect 442 182 447 189
rect 453 187 460 189
rect 453 185 455 187
rect 457 185 460 187
rect 442 180 449 182
rect 442 178 445 180
rect 447 178 449 180
rect 442 176 449 178
rect 453 180 460 185
rect 453 178 455 180
rect 457 178 460 180
rect 442 169 447 176
rect 453 175 460 178
rect 462 187 470 189
rect 462 185 465 187
rect 467 185 470 187
rect 462 175 470 185
rect 472 182 477 189
rect 527 183 534 189
rect 472 179 480 182
rect 472 177 475 179
rect 477 177 480 179
rect 472 175 480 177
rect 475 172 480 175
rect 482 176 490 182
rect 482 174 485 176
rect 487 174 490 176
rect 482 172 490 174
rect 485 169 490 172
rect 492 180 499 182
rect 492 178 495 180
rect 497 178 499 180
rect 492 176 499 178
rect 516 180 523 183
rect 516 178 518 180
rect 520 178 523 180
rect 516 176 523 178
rect 492 169 497 176
rect 518 169 523 176
rect 525 173 534 183
rect 525 171 529 173
rect 531 171 534 173
rect 525 169 534 171
rect 536 169 541 189
rect 543 182 548 189
rect 554 187 561 189
rect 554 185 556 187
rect 558 185 561 187
rect 543 180 550 182
rect 543 178 546 180
rect 548 178 550 180
rect 543 176 550 178
rect 554 180 561 185
rect 554 178 556 180
rect 558 178 561 180
rect 543 169 548 176
rect 554 175 561 178
rect 563 187 571 189
rect 563 185 566 187
rect 568 185 571 187
rect 563 175 571 185
rect 573 182 578 189
rect 626 183 633 189
rect 573 179 581 182
rect 573 177 576 179
rect 578 177 581 179
rect 573 175 581 177
rect 576 172 581 175
rect 583 176 591 182
rect 583 174 586 176
rect 588 174 591 176
rect 583 172 591 174
rect 586 169 591 172
rect 593 180 600 182
rect 593 178 596 180
rect 598 178 600 180
rect 593 176 600 178
rect 615 180 622 183
rect 615 178 617 180
rect 619 178 622 180
rect 615 176 622 178
rect 593 169 598 176
rect 617 169 622 176
rect 624 173 633 183
rect 624 171 628 173
rect 630 171 633 173
rect 624 169 633 171
rect 635 169 640 189
rect 642 182 647 189
rect 653 187 660 189
rect 653 185 655 187
rect 657 185 660 187
rect 642 180 649 182
rect 642 178 645 180
rect 647 178 649 180
rect 642 176 649 178
rect 653 180 660 185
rect 653 178 655 180
rect 657 178 660 180
rect 642 169 647 176
rect 653 175 660 178
rect 662 187 670 189
rect 662 185 665 187
rect 667 185 670 187
rect 662 175 670 185
rect 672 182 677 189
rect 672 179 680 182
rect 672 177 675 179
rect 677 177 680 179
rect 672 175 680 177
rect 675 172 680 175
rect 682 176 690 182
rect 682 174 685 176
rect 687 174 690 176
rect 682 172 690 174
rect 685 169 690 172
rect 692 180 699 182
rect 692 178 695 180
rect 697 178 699 180
rect 692 176 699 178
rect 692 169 697 176
rect 22 150 27 157
rect 20 148 27 150
rect 20 146 22 148
rect 24 146 27 148
rect 20 143 27 146
rect 29 155 38 157
rect 29 153 33 155
rect 35 153 38 155
rect 29 143 38 153
rect 31 137 38 143
rect 40 137 45 157
rect 47 150 52 157
rect 90 154 95 157
rect 80 151 85 154
rect 47 148 54 150
rect 47 146 50 148
rect 52 146 54 148
rect 47 144 54 146
rect 58 148 65 151
rect 58 146 60 148
rect 62 146 65 148
rect 47 137 52 144
rect 58 141 65 146
rect 58 139 60 141
rect 62 139 65 141
rect 58 137 65 139
rect 67 141 75 151
rect 67 139 70 141
rect 72 139 75 141
rect 67 137 75 139
rect 77 149 85 151
rect 77 147 80 149
rect 82 147 85 149
rect 77 144 85 147
rect 87 152 95 154
rect 87 150 90 152
rect 92 150 95 152
rect 87 144 95 150
rect 97 150 102 157
rect 97 148 104 150
rect 97 146 100 148
rect 102 146 104 148
rect 97 144 104 146
rect 108 148 115 151
rect 108 146 110 148
rect 112 146 115 148
rect 77 137 82 144
rect 108 141 115 146
rect 108 139 110 141
rect 112 139 115 141
rect 108 137 115 139
rect 117 150 122 151
rect 117 148 125 150
rect 117 146 120 148
rect 122 146 125 148
rect 117 142 125 146
rect 127 148 132 150
rect 163 150 168 157
rect 161 148 168 150
rect 127 146 135 148
rect 127 144 130 146
rect 132 144 135 146
rect 127 142 135 144
rect 117 137 122 142
rect 130 140 135 142
rect 137 146 144 148
rect 137 144 140 146
rect 142 144 144 146
rect 137 140 144 144
rect 161 146 163 148
rect 165 146 168 148
rect 161 143 168 146
rect 170 155 179 157
rect 170 153 174 155
rect 176 153 179 155
rect 170 143 179 153
rect 172 137 179 143
rect 181 137 186 157
rect 188 150 193 157
rect 231 154 236 157
rect 221 151 226 154
rect 188 148 195 150
rect 188 146 191 148
rect 193 146 195 148
rect 188 144 195 146
rect 199 148 206 151
rect 199 146 201 148
rect 203 146 206 148
rect 188 137 193 144
rect 199 141 206 146
rect 199 139 201 141
rect 203 139 206 141
rect 199 137 206 139
rect 208 141 216 151
rect 208 139 211 141
rect 213 139 216 141
rect 208 137 216 139
rect 218 149 226 151
rect 218 147 221 149
rect 223 147 226 149
rect 218 144 226 147
rect 228 152 236 154
rect 228 150 231 152
rect 233 150 236 152
rect 228 144 236 150
rect 238 150 243 157
rect 263 150 268 157
rect 238 148 245 150
rect 238 146 241 148
rect 243 146 245 148
rect 238 144 245 146
rect 261 148 268 150
rect 261 146 263 148
rect 265 146 268 148
rect 261 144 268 146
rect 270 154 275 157
rect 270 152 278 154
rect 270 150 273 152
rect 275 150 278 152
rect 270 144 278 150
rect 280 151 285 154
rect 280 149 288 151
rect 280 147 283 149
rect 285 147 288 149
rect 280 144 288 147
rect 218 137 223 144
rect 283 137 288 144
rect 290 141 298 151
rect 290 139 293 141
rect 295 139 298 141
rect 290 137 298 139
rect 300 148 307 151
rect 313 150 318 157
rect 300 146 303 148
rect 305 146 307 148
rect 300 141 307 146
rect 311 148 318 150
rect 311 146 313 148
rect 315 146 318 148
rect 311 144 318 146
rect 300 139 303 141
rect 305 139 307 141
rect 300 137 307 139
rect 313 137 318 144
rect 320 137 325 157
rect 327 155 336 157
rect 327 153 330 155
rect 332 153 336 155
rect 327 143 336 153
rect 338 150 343 157
rect 338 148 345 150
rect 338 146 341 148
rect 343 146 345 148
rect 338 143 345 146
rect 362 148 369 151
rect 362 146 364 148
rect 366 146 369 148
rect 327 137 334 143
rect 362 141 369 146
rect 362 139 364 141
rect 366 139 369 141
rect 362 137 369 139
rect 371 150 376 151
rect 371 148 379 150
rect 371 146 374 148
rect 376 146 379 148
rect 371 142 379 146
rect 381 148 386 150
rect 417 150 422 157
rect 415 148 422 150
rect 381 146 389 148
rect 381 144 384 146
rect 386 144 389 146
rect 381 142 389 144
rect 371 137 376 142
rect 384 140 389 142
rect 391 146 398 148
rect 391 144 394 146
rect 396 144 398 146
rect 391 140 398 144
rect 415 146 417 148
rect 419 146 422 148
rect 415 143 422 146
rect 424 155 433 157
rect 424 153 428 155
rect 430 153 433 155
rect 424 143 433 153
rect 426 137 433 143
rect 435 137 440 157
rect 442 150 447 157
rect 485 154 490 157
rect 475 151 480 154
rect 442 148 449 150
rect 442 146 445 148
rect 447 146 449 148
rect 442 144 449 146
rect 453 148 460 151
rect 453 146 455 148
rect 457 146 460 148
rect 442 137 447 144
rect 453 141 460 146
rect 453 139 455 141
rect 457 139 460 141
rect 453 137 460 139
rect 462 141 470 151
rect 462 139 465 141
rect 467 139 470 141
rect 462 137 470 139
rect 472 149 480 151
rect 472 147 475 149
rect 477 147 480 149
rect 472 144 480 147
rect 482 152 490 154
rect 482 150 485 152
rect 487 150 490 152
rect 482 144 490 150
rect 492 150 497 157
rect 518 150 523 157
rect 492 148 499 150
rect 492 146 495 148
rect 497 146 499 148
rect 492 144 499 146
rect 516 148 523 150
rect 516 146 518 148
rect 520 146 523 148
rect 472 137 477 144
rect 516 143 523 146
rect 525 155 534 157
rect 525 153 529 155
rect 531 153 534 155
rect 525 143 534 153
rect 527 137 534 143
rect 536 137 541 157
rect 543 150 548 157
rect 586 154 591 157
rect 576 151 581 154
rect 543 148 550 150
rect 543 146 546 148
rect 548 146 550 148
rect 543 144 550 146
rect 554 148 561 151
rect 554 146 556 148
rect 558 146 561 148
rect 543 137 548 144
rect 554 141 561 146
rect 554 139 556 141
rect 558 139 561 141
rect 554 137 561 139
rect 563 141 571 151
rect 563 139 566 141
rect 568 139 571 141
rect 563 137 571 139
rect 573 149 581 151
rect 573 147 576 149
rect 578 147 581 149
rect 573 144 581 147
rect 583 152 591 154
rect 583 150 586 152
rect 588 150 591 152
rect 583 144 591 150
rect 593 150 598 157
rect 617 150 622 157
rect 593 148 600 150
rect 593 146 596 148
rect 598 146 600 148
rect 593 144 600 146
rect 615 148 622 150
rect 615 146 617 148
rect 619 146 622 148
rect 573 137 578 144
rect 615 143 622 146
rect 624 155 633 157
rect 624 153 628 155
rect 630 153 633 155
rect 624 143 633 153
rect 626 137 633 143
rect 635 137 640 157
rect 642 150 647 157
rect 685 154 690 157
rect 675 151 680 154
rect 642 148 649 150
rect 642 146 645 148
rect 647 146 649 148
rect 642 144 649 146
rect 653 148 660 151
rect 653 146 655 148
rect 657 146 660 148
rect 642 137 647 144
rect 653 141 660 146
rect 653 139 655 141
rect 657 139 660 141
rect 653 137 660 139
rect 662 141 670 151
rect 662 139 665 141
rect 667 139 670 141
rect 662 137 670 139
rect 672 149 680 151
rect 672 147 675 149
rect 677 147 680 149
rect 672 144 680 147
rect 682 152 690 154
rect 682 150 685 152
rect 687 150 690 152
rect 682 144 690 150
rect 692 150 697 157
rect 692 148 699 150
rect 692 146 695 148
rect 697 146 699 148
rect 692 144 699 146
rect 672 137 677 144
rect 18 43 25 45
rect 18 41 20 43
rect 22 41 25 43
rect 18 36 25 41
rect 18 34 20 36
rect 22 34 25 36
rect 18 31 25 34
rect 27 40 32 45
rect 40 40 45 42
rect 27 36 35 40
rect 27 34 30 36
rect 32 34 35 36
rect 27 32 35 34
rect 37 38 45 40
rect 37 36 40 38
rect 42 36 45 38
rect 37 34 45 36
rect 47 38 54 42
rect 70 39 77 45
rect 47 36 50 38
rect 52 36 54 38
rect 47 34 54 36
rect 59 36 66 39
rect 59 34 61 36
rect 63 34 66 36
rect 37 32 42 34
rect 27 31 32 32
rect 59 32 66 34
rect 61 25 66 32
rect 68 29 77 39
rect 68 27 72 29
rect 74 27 77 29
rect 68 25 77 27
rect 79 25 84 45
rect 86 38 91 45
rect 97 43 104 45
rect 97 41 99 43
rect 101 41 104 43
rect 86 36 93 38
rect 86 34 89 36
rect 91 34 93 36
rect 86 32 93 34
rect 97 36 104 41
rect 97 34 99 36
rect 101 34 104 36
rect 86 25 91 32
rect 97 31 104 34
rect 106 43 114 45
rect 106 41 109 43
rect 111 41 114 43
rect 106 31 114 41
rect 116 38 121 45
rect 171 39 178 45
rect 116 35 124 38
rect 116 33 119 35
rect 121 33 124 35
rect 116 31 124 33
rect 119 28 124 31
rect 126 32 134 38
rect 126 30 129 32
rect 131 30 134 32
rect 126 28 134 30
rect 129 25 134 28
rect 136 36 143 38
rect 136 34 139 36
rect 141 34 143 36
rect 136 32 143 34
rect 160 36 167 39
rect 160 34 162 36
rect 164 34 167 36
rect 160 32 167 34
rect 136 25 141 32
rect 162 25 167 32
rect 169 29 178 39
rect 169 27 173 29
rect 175 27 178 29
rect 169 25 178 27
rect 180 25 185 45
rect 187 38 192 45
rect 198 43 205 45
rect 198 41 200 43
rect 202 41 205 43
rect 187 36 194 38
rect 187 34 190 36
rect 192 34 194 36
rect 187 32 194 34
rect 198 36 205 41
rect 198 34 200 36
rect 202 34 205 36
rect 187 25 192 32
rect 198 31 205 34
rect 207 43 215 45
rect 207 41 210 43
rect 212 41 215 43
rect 207 31 215 41
rect 217 38 222 45
rect 272 39 279 45
rect 217 35 225 38
rect 217 33 220 35
rect 222 33 225 35
rect 217 31 225 33
rect 220 28 225 31
rect 227 32 235 38
rect 227 30 230 32
rect 232 30 235 32
rect 227 28 235 30
rect 230 25 235 28
rect 237 36 244 38
rect 237 34 240 36
rect 242 34 244 36
rect 237 32 244 34
rect 261 36 268 39
rect 261 34 263 36
rect 265 34 268 36
rect 261 32 268 34
rect 237 25 242 32
rect 263 25 268 32
rect 270 29 279 39
rect 270 27 274 29
rect 276 27 279 29
rect 270 25 279 27
rect 281 25 286 45
rect 288 38 293 45
rect 299 43 306 45
rect 299 41 301 43
rect 303 41 306 43
rect 288 36 295 38
rect 288 34 291 36
rect 293 34 295 36
rect 288 32 295 34
rect 299 36 306 41
rect 299 34 301 36
rect 303 34 306 36
rect 288 25 293 32
rect 299 31 306 34
rect 308 43 316 45
rect 308 41 311 43
rect 313 41 316 43
rect 308 31 316 41
rect 318 38 323 45
rect 361 43 368 45
rect 361 41 363 43
rect 365 41 368 43
rect 318 35 326 38
rect 318 33 321 35
rect 323 33 326 35
rect 318 31 326 33
rect 321 28 326 31
rect 328 32 336 38
rect 328 30 331 32
rect 333 30 336 32
rect 328 28 336 30
rect 331 25 336 28
rect 338 36 345 38
rect 338 34 341 36
rect 343 34 345 36
rect 338 32 345 34
rect 361 36 368 41
rect 361 34 363 36
rect 365 34 368 36
rect 338 25 343 32
rect 361 31 368 34
rect 370 40 375 45
rect 383 40 388 42
rect 370 36 378 40
rect 370 34 373 36
rect 375 34 378 36
rect 370 32 378 34
rect 380 38 388 40
rect 380 36 383 38
rect 385 36 388 38
rect 380 34 388 36
rect 390 38 397 42
rect 425 39 432 45
rect 390 36 393 38
rect 395 36 397 38
rect 390 34 397 36
rect 414 36 421 39
rect 414 34 416 36
rect 418 34 421 36
rect 380 32 385 34
rect 370 31 375 32
rect 414 32 421 34
rect 416 25 421 32
rect 423 29 432 39
rect 423 27 427 29
rect 429 27 432 29
rect 423 25 432 27
rect 434 25 439 45
rect 441 38 446 45
rect 452 43 459 45
rect 452 41 454 43
rect 456 41 459 43
rect 441 36 448 38
rect 441 34 444 36
rect 446 34 448 36
rect 441 32 448 34
rect 452 36 459 41
rect 452 34 454 36
rect 456 34 459 36
rect 441 25 446 32
rect 452 31 459 34
rect 461 43 469 45
rect 461 41 464 43
rect 466 41 469 43
rect 461 31 469 41
rect 471 38 476 45
rect 526 39 533 45
rect 471 35 479 38
rect 471 33 474 35
rect 476 33 479 35
rect 471 31 479 33
rect 474 28 479 31
rect 481 32 489 38
rect 481 30 484 32
rect 486 30 489 32
rect 481 28 489 30
rect 484 25 489 28
rect 491 36 498 38
rect 491 34 494 36
rect 496 34 498 36
rect 491 32 498 34
rect 515 36 522 39
rect 515 34 517 36
rect 519 34 522 36
rect 515 32 522 34
rect 491 25 496 32
rect 517 25 522 32
rect 524 29 533 39
rect 524 27 528 29
rect 530 27 533 29
rect 524 25 533 27
rect 535 25 540 45
rect 542 38 547 45
rect 553 43 560 45
rect 553 41 555 43
rect 557 41 560 43
rect 542 36 549 38
rect 542 34 545 36
rect 547 34 549 36
rect 542 32 549 34
rect 553 36 560 41
rect 553 34 555 36
rect 557 34 560 36
rect 542 25 547 32
rect 553 31 560 34
rect 562 43 570 45
rect 562 41 565 43
rect 567 41 570 43
rect 562 31 570 41
rect 572 38 577 45
rect 625 39 632 45
rect 572 35 580 38
rect 572 33 575 35
rect 577 33 580 35
rect 572 31 580 33
rect 575 28 580 31
rect 582 32 590 38
rect 582 30 585 32
rect 587 30 590 32
rect 582 28 590 30
rect 585 25 590 28
rect 592 36 599 38
rect 592 34 595 36
rect 597 34 599 36
rect 592 32 599 34
rect 614 36 621 39
rect 614 34 616 36
rect 618 34 621 36
rect 614 32 621 34
rect 592 25 597 32
rect 616 25 621 32
rect 623 29 632 39
rect 623 27 627 29
rect 629 27 632 29
rect 623 25 632 27
rect 634 25 639 45
rect 641 38 646 45
rect 652 43 659 45
rect 652 41 654 43
rect 656 41 659 43
rect 641 36 648 38
rect 641 34 644 36
rect 646 34 648 36
rect 641 32 648 34
rect 652 36 659 41
rect 652 34 654 36
rect 656 34 659 36
rect 641 25 646 32
rect 652 31 659 34
rect 661 43 669 45
rect 661 41 664 43
rect 666 41 669 43
rect 661 31 669 41
rect 671 38 676 45
rect 671 35 679 38
rect 671 33 674 35
rect 676 33 679 35
rect 671 31 679 33
rect 674 28 679 31
rect 681 32 689 38
rect 681 30 684 32
rect 686 30 689 32
rect 681 28 689 30
rect 684 25 689 28
rect 691 36 698 38
rect 691 34 694 36
rect 696 34 698 36
rect 691 32 698 34
rect 691 25 696 32
<< pdif >>
rect 18 371 25 373
rect 18 369 20 371
rect 22 369 25 371
rect 18 364 25 369
rect 18 362 20 364
rect 22 362 25 364
rect 18 354 25 362
rect 27 365 35 373
rect 27 363 30 365
rect 32 363 35 365
rect 27 358 35 363
rect 27 356 30 358
rect 32 356 35 358
rect 27 354 35 356
rect 37 371 45 373
rect 37 369 40 371
rect 42 369 45 371
rect 37 364 45 369
rect 37 362 40 364
rect 42 362 45 364
rect 37 354 45 362
rect 39 345 45 354
rect 47 366 52 373
rect 58 371 65 373
rect 58 369 60 371
rect 62 369 65 371
rect 47 364 54 366
rect 47 362 50 364
rect 52 362 54 364
rect 47 357 54 362
rect 47 355 50 357
rect 52 355 54 357
rect 47 353 54 355
rect 58 364 65 369
rect 58 362 60 364
rect 62 362 65 364
rect 58 354 65 362
rect 67 365 75 373
rect 67 363 70 365
rect 72 363 75 365
rect 67 358 75 363
rect 67 356 70 358
rect 72 356 75 358
rect 67 354 75 356
rect 77 371 85 373
rect 77 369 80 371
rect 82 369 85 371
rect 77 364 85 369
rect 77 362 80 364
rect 82 362 85 364
rect 77 354 85 362
rect 47 345 52 353
rect 79 345 85 354
rect 87 366 92 373
rect 87 364 94 366
rect 87 362 90 364
rect 92 362 94 364
rect 87 357 94 362
rect 101 358 106 373
rect 87 355 90 357
rect 92 355 94 357
rect 87 353 94 355
rect 99 356 106 358
rect 99 354 101 356
rect 103 354 106 356
rect 87 345 92 353
rect 99 349 106 354
rect 99 347 101 349
rect 103 347 106 349
rect 99 345 106 347
rect 108 371 116 373
rect 108 369 111 371
rect 113 369 116 371
rect 108 364 116 369
rect 108 362 111 364
rect 113 362 116 364
rect 108 345 116 362
rect 118 363 126 373
rect 118 361 121 363
rect 123 361 126 363
rect 118 356 126 361
rect 118 354 121 356
rect 123 354 126 356
rect 118 345 126 354
rect 128 371 142 373
rect 128 369 133 371
rect 135 370 142 371
rect 165 371 174 373
rect 135 369 144 370
rect 128 364 144 369
rect 128 362 133 364
rect 135 362 144 364
rect 128 345 144 362
rect 146 345 151 370
rect 153 361 158 370
rect 165 369 168 371
rect 170 369 174 371
rect 165 361 174 369
rect 153 352 161 361
rect 153 350 156 352
rect 158 350 161 352
rect 153 348 161 350
rect 163 348 174 361
rect 176 361 181 373
rect 197 361 202 373
rect 176 359 183 361
rect 176 357 179 359
rect 181 357 183 359
rect 176 352 183 357
rect 176 350 179 352
rect 181 350 183 352
rect 176 348 183 350
rect 195 359 202 361
rect 195 357 197 359
rect 199 357 202 359
rect 195 352 202 357
rect 195 350 197 352
rect 199 350 202 352
rect 195 348 202 350
rect 204 371 213 373
rect 204 369 208 371
rect 210 369 213 371
rect 236 371 250 373
rect 236 370 243 371
rect 204 361 213 369
rect 220 361 225 370
rect 204 348 215 361
rect 217 352 225 361
rect 217 350 220 352
rect 222 350 225 352
rect 217 348 225 350
rect 153 345 158 348
rect 220 345 225 348
rect 227 345 232 370
rect 234 369 243 370
rect 245 369 250 371
rect 234 364 250 369
rect 234 362 243 364
rect 245 362 250 364
rect 234 345 250 362
rect 252 363 260 373
rect 252 361 255 363
rect 257 361 260 363
rect 252 356 260 361
rect 252 354 255 356
rect 257 354 260 356
rect 252 345 260 354
rect 262 371 270 373
rect 262 369 265 371
rect 267 369 270 371
rect 262 364 270 369
rect 262 362 265 364
rect 267 362 270 364
rect 262 345 270 362
rect 272 358 277 373
rect 286 366 291 373
rect 284 364 291 366
rect 284 362 286 364
rect 288 362 291 364
rect 272 356 279 358
rect 272 354 275 356
rect 277 354 279 356
rect 272 349 279 354
rect 284 357 291 362
rect 284 355 286 357
rect 288 355 291 357
rect 284 353 291 355
rect 272 347 275 349
rect 277 347 279 349
rect 272 345 279 347
rect 286 345 291 353
rect 293 371 301 373
rect 293 369 296 371
rect 298 369 301 371
rect 293 364 301 369
rect 293 362 296 364
rect 298 362 301 364
rect 293 354 301 362
rect 303 365 311 373
rect 303 363 306 365
rect 308 363 311 365
rect 303 358 311 363
rect 303 356 306 358
rect 308 356 311 358
rect 303 354 311 356
rect 313 371 320 373
rect 313 369 316 371
rect 318 369 320 371
rect 313 364 320 369
rect 326 366 331 373
rect 313 362 316 364
rect 318 362 320 364
rect 313 354 320 362
rect 324 364 331 366
rect 324 362 326 364
rect 328 362 331 364
rect 324 357 331 362
rect 324 355 326 357
rect 328 355 331 357
rect 293 345 299 354
rect 324 353 331 355
rect 326 345 331 353
rect 333 371 341 373
rect 333 369 336 371
rect 338 369 341 371
rect 333 364 341 369
rect 333 362 336 364
rect 338 362 341 364
rect 333 354 341 362
rect 343 365 351 373
rect 343 363 346 365
rect 348 363 351 365
rect 343 358 351 363
rect 343 356 346 358
rect 348 356 351 358
rect 343 354 351 356
rect 353 371 360 373
rect 353 369 356 371
rect 358 369 360 371
rect 353 364 360 369
rect 353 362 356 364
rect 358 362 360 364
rect 353 354 360 362
rect 367 361 372 373
rect 365 359 372 361
rect 365 357 367 359
rect 369 357 372 359
rect 333 345 339 354
rect 365 352 372 357
rect 365 350 367 352
rect 369 350 372 352
rect 365 348 372 350
rect 374 371 383 373
rect 374 369 378 371
rect 380 369 383 371
rect 406 371 420 373
rect 406 370 413 371
rect 374 361 383 369
rect 390 361 395 370
rect 374 348 385 361
rect 387 352 395 361
rect 387 350 390 352
rect 392 350 395 352
rect 387 348 395 350
rect 390 345 395 348
rect 397 345 402 370
rect 404 369 413 370
rect 415 369 420 371
rect 404 364 420 369
rect 404 362 413 364
rect 415 362 420 364
rect 404 345 420 362
rect 422 363 430 373
rect 422 361 425 363
rect 427 361 430 363
rect 422 356 430 361
rect 422 354 425 356
rect 427 354 430 356
rect 422 345 430 354
rect 432 371 440 373
rect 432 369 435 371
rect 437 369 440 371
rect 432 364 440 369
rect 432 362 435 364
rect 437 362 440 364
rect 432 345 440 362
rect 442 358 447 373
rect 456 366 461 373
rect 454 364 461 366
rect 454 362 456 364
rect 458 362 461 364
rect 442 356 449 358
rect 442 354 445 356
rect 447 354 449 356
rect 442 349 449 354
rect 454 357 461 362
rect 454 355 456 357
rect 458 355 461 357
rect 454 353 461 355
rect 442 347 445 349
rect 447 347 449 349
rect 442 345 449 347
rect 456 345 461 353
rect 463 371 471 373
rect 463 369 466 371
rect 468 369 471 371
rect 463 364 471 369
rect 463 362 466 364
rect 468 362 471 364
rect 463 354 471 362
rect 473 365 481 373
rect 473 363 476 365
rect 478 363 481 365
rect 473 358 481 363
rect 473 356 476 358
rect 478 356 481 358
rect 473 354 481 356
rect 483 371 490 373
rect 483 369 486 371
rect 488 369 490 371
rect 483 364 490 369
rect 496 366 501 373
rect 483 362 486 364
rect 488 362 490 364
rect 483 354 490 362
rect 494 364 501 366
rect 494 362 496 364
rect 498 362 501 364
rect 494 357 501 362
rect 494 355 496 357
rect 498 355 501 357
rect 463 345 469 354
rect 494 353 501 355
rect 496 345 501 353
rect 503 371 511 373
rect 503 369 506 371
rect 508 369 511 371
rect 503 364 511 369
rect 503 362 506 364
rect 508 362 511 364
rect 503 354 511 362
rect 513 365 521 373
rect 513 363 516 365
rect 518 363 521 365
rect 513 358 521 363
rect 513 356 516 358
rect 518 356 521 358
rect 513 354 521 356
rect 523 371 530 373
rect 523 369 526 371
rect 528 369 530 371
rect 523 364 530 369
rect 523 362 526 364
rect 528 362 530 364
rect 523 354 530 362
rect 534 371 541 373
rect 534 369 536 371
rect 538 369 541 371
rect 534 364 541 369
rect 534 362 536 364
rect 538 362 541 364
rect 534 354 541 362
rect 543 365 551 373
rect 543 363 546 365
rect 548 363 551 365
rect 543 358 551 363
rect 543 356 546 358
rect 548 356 551 358
rect 543 354 551 356
rect 553 371 561 373
rect 553 369 556 371
rect 558 369 561 371
rect 553 364 561 369
rect 553 362 556 364
rect 558 362 561 364
rect 553 354 561 362
rect 503 345 509 354
rect 555 345 561 354
rect 563 366 568 373
rect 574 371 581 373
rect 574 369 576 371
rect 578 369 581 371
rect 563 364 570 366
rect 563 362 566 364
rect 568 362 570 364
rect 563 357 570 362
rect 563 355 566 357
rect 568 355 570 357
rect 563 353 570 355
rect 574 364 581 369
rect 574 362 576 364
rect 578 362 581 364
rect 574 354 581 362
rect 583 365 591 373
rect 583 363 586 365
rect 588 363 591 365
rect 583 358 591 363
rect 583 356 586 358
rect 588 356 591 358
rect 583 354 591 356
rect 593 371 601 373
rect 593 369 596 371
rect 598 369 601 371
rect 593 364 601 369
rect 593 362 596 364
rect 598 362 601 364
rect 593 354 601 362
rect 563 345 568 353
rect 595 345 601 354
rect 603 366 608 373
rect 603 364 610 366
rect 603 362 606 364
rect 608 362 610 364
rect 603 357 610 362
rect 617 358 622 373
rect 603 355 606 357
rect 608 355 610 357
rect 603 353 610 355
rect 615 356 622 358
rect 615 354 617 356
rect 619 354 622 356
rect 603 345 608 353
rect 615 349 622 354
rect 615 347 617 349
rect 619 347 622 349
rect 615 345 622 347
rect 624 371 632 373
rect 624 369 627 371
rect 629 369 632 371
rect 624 364 632 369
rect 624 362 627 364
rect 629 362 632 364
rect 624 345 632 362
rect 634 363 642 373
rect 634 361 637 363
rect 639 361 642 363
rect 634 356 642 361
rect 634 354 637 356
rect 639 354 642 356
rect 634 345 642 354
rect 644 371 658 373
rect 644 369 649 371
rect 651 370 658 371
rect 681 371 690 373
rect 651 369 660 370
rect 644 364 660 369
rect 644 362 649 364
rect 651 362 660 364
rect 644 345 660 362
rect 662 345 667 370
rect 669 361 674 370
rect 681 369 684 371
rect 686 369 690 371
rect 681 361 690 369
rect 669 352 677 361
rect 669 350 672 352
rect 674 350 677 352
rect 669 348 677 350
rect 679 348 690 361
rect 692 361 697 373
rect 692 359 699 361
rect 692 357 695 359
rect 697 357 699 359
rect 692 352 699 357
rect 692 350 695 352
rect 697 350 699 352
rect 692 348 699 350
rect 669 345 674 348
rect 39 260 45 269
rect 18 252 25 260
rect 18 250 20 252
rect 22 250 25 252
rect 18 245 25 250
rect 18 243 20 245
rect 22 243 25 245
rect 18 241 25 243
rect 27 258 35 260
rect 27 256 30 258
rect 32 256 35 258
rect 27 251 35 256
rect 27 249 30 251
rect 32 249 35 251
rect 27 241 35 249
rect 37 252 45 260
rect 37 250 40 252
rect 42 250 45 252
rect 37 245 45 250
rect 37 243 40 245
rect 42 243 45 245
rect 37 241 45 243
rect 47 261 52 269
rect 47 259 54 261
rect 79 260 85 269
rect 47 257 50 259
rect 52 257 54 259
rect 47 252 54 257
rect 47 250 50 252
rect 52 250 54 252
rect 47 248 54 250
rect 58 252 65 260
rect 58 250 60 252
rect 62 250 65 252
rect 47 241 52 248
rect 58 245 65 250
rect 58 243 60 245
rect 62 243 65 245
rect 58 241 65 243
rect 67 258 75 260
rect 67 256 70 258
rect 72 256 75 258
rect 67 251 75 256
rect 67 249 70 251
rect 72 249 75 251
rect 67 241 75 249
rect 77 252 85 260
rect 77 250 80 252
rect 82 250 85 252
rect 77 245 85 250
rect 77 243 80 245
rect 82 243 85 245
rect 77 241 85 243
rect 87 261 92 269
rect 99 267 106 269
rect 99 265 101 267
rect 103 265 106 267
rect 87 259 94 261
rect 87 257 90 259
rect 92 257 94 259
rect 87 252 94 257
rect 99 256 106 265
rect 87 250 90 252
rect 92 250 94 252
rect 87 248 94 250
rect 87 241 92 248
rect 101 241 106 256
rect 108 252 116 269
rect 108 250 111 252
rect 113 250 116 252
rect 108 245 116 250
rect 108 243 111 245
rect 113 243 116 245
rect 108 241 116 243
rect 118 260 126 269
rect 118 258 121 260
rect 123 258 126 260
rect 118 253 126 258
rect 118 251 121 253
rect 123 251 126 253
rect 118 241 126 251
rect 128 252 144 269
rect 128 250 133 252
rect 135 250 144 252
rect 128 245 144 250
rect 128 243 133 245
rect 135 244 144 245
rect 146 244 151 269
rect 153 266 158 269
rect 220 266 225 269
rect 153 264 161 266
rect 153 262 156 264
rect 158 262 161 264
rect 153 253 161 262
rect 163 253 174 266
rect 153 244 158 253
rect 165 245 174 253
rect 135 243 142 244
rect 128 241 142 243
rect 165 243 168 245
rect 170 243 174 245
rect 165 241 174 243
rect 176 264 183 266
rect 176 262 179 264
rect 181 262 183 264
rect 176 257 183 262
rect 176 255 179 257
rect 181 255 183 257
rect 176 253 183 255
rect 195 264 202 266
rect 195 262 197 264
rect 199 262 202 264
rect 195 257 202 262
rect 195 255 197 257
rect 199 255 202 257
rect 195 253 202 255
rect 176 241 181 253
rect 197 241 202 253
rect 204 253 215 266
rect 217 264 225 266
rect 217 262 220 264
rect 222 262 225 264
rect 217 253 225 262
rect 204 245 213 253
rect 204 243 208 245
rect 210 243 213 245
rect 220 244 225 253
rect 227 244 232 269
rect 234 252 250 269
rect 234 250 243 252
rect 245 250 250 252
rect 234 245 250 250
rect 234 244 243 245
rect 204 241 213 243
rect 236 243 243 244
rect 245 243 250 245
rect 236 241 250 243
rect 252 260 260 269
rect 252 258 255 260
rect 257 258 260 260
rect 252 253 260 258
rect 252 251 255 253
rect 257 251 260 253
rect 252 241 260 251
rect 262 252 270 269
rect 262 250 265 252
rect 267 250 270 252
rect 262 245 270 250
rect 262 243 265 245
rect 267 243 270 245
rect 262 241 270 243
rect 272 267 279 269
rect 272 265 275 267
rect 277 265 279 267
rect 272 260 279 265
rect 286 261 291 269
rect 272 258 275 260
rect 277 258 279 260
rect 272 256 279 258
rect 284 259 291 261
rect 284 257 286 259
rect 288 257 291 259
rect 272 241 277 256
rect 284 252 291 257
rect 284 250 286 252
rect 288 250 291 252
rect 284 248 291 250
rect 286 241 291 248
rect 293 260 299 269
rect 326 261 331 269
rect 293 252 301 260
rect 293 250 296 252
rect 298 250 301 252
rect 293 245 301 250
rect 293 243 296 245
rect 298 243 301 245
rect 293 241 301 243
rect 303 258 311 260
rect 303 256 306 258
rect 308 256 311 258
rect 303 251 311 256
rect 303 249 306 251
rect 308 249 311 251
rect 303 241 311 249
rect 313 252 320 260
rect 313 250 316 252
rect 318 250 320 252
rect 313 245 320 250
rect 324 259 331 261
rect 324 257 326 259
rect 328 257 331 259
rect 324 252 331 257
rect 324 250 326 252
rect 328 250 331 252
rect 324 248 331 250
rect 313 243 316 245
rect 318 243 320 245
rect 313 241 320 243
rect 326 241 331 248
rect 333 260 339 269
rect 390 266 395 269
rect 365 264 372 266
rect 365 262 367 264
rect 369 262 372 264
rect 333 252 341 260
rect 333 250 336 252
rect 338 250 341 252
rect 333 245 341 250
rect 333 243 336 245
rect 338 243 341 245
rect 333 241 341 243
rect 343 258 351 260
rect 343 256 346 258
rect 348 256 351 258
rect 343 251 351 256
rect 343 249 346 251
rect 348 249 351 251
rect 343 241 351 249
rect 353 252 360 260
rect 365 257 372 262
rect 365 255 367 257
rect 369 255 372 257
rect 365 253 372 255
rect 353 250 356 252
rect 358 250 360 252
rect 353 245 360 250
rect 353 243 356 245
rect 358 243 360 245
rect 353 241 360 243
rect 367 241 372 253
rect 374 253 385 266
rect 387 264 395 266
rect 387 262 390 264
rect 392 262 395 264
rect 387 253 395 262
rect 374 245 383 253
rect 374 243 378 245
rect 380 243 383 245
rect 390 244 395 253
rect 397 244 402 269
rect 404 252 420 269
rect 404 250 413 252
rect 415 250 420 252
rect 404 245 420 250
rect 404 244 413 245
rect 374 241 383 243
rect 406 243 413 244
rect 415 243 420 245
rect 406 241 420 243
rect 422 260 430 269
rect 422 258 425 260
rect 427 258 430 260
rect 422 253 430 258
rect 422 251 425 253
rect 427 251 430 253
rect 422 241 430 251
rect 432 252 440 269
rect 432 250 435 252
rect 437 250 440 252
rect 432 245 440 250
rect 432 243 435 245
rect 437 243 440 245
rect 432 241 440 243
rect 442 267 449 269
rect 442 265 445 267
rect 447 265 449 267
rect 442 260 449 265
rect 456 261 461 269
rect 442 258 445 260
rect 447 258 449 260
rect 442 256 449 258
rect 454 259 461 261
rect 454 257 456 259
rect 458 257 461 259
rect 442 241 447 256
rect 454 252 461 257
rect 454 250 456 252
rect 458 250 461 252
rect 454 248 461 250
rect 456 241 461 248
rect 463 260 469 269
rect 496 261 501 269
rect 463 252 471 260
rect 463 250 466 252
rect 468 250 471 252
rect 463 245 471 250
rect 463 243 466 245
rect 468 243 471 245
rect 463 241 471 243
rect 473 258 481 260
rect 473 256 476 258
rect 478 256 481 258
rect 473 251 481 256
rect 473 249 476 251
rect 478 249 481 251
rect 473 241 481 249
rect 483 252 490 260
rect 483 250 486 252
rect 488 250 490 252
rect 483 245 490 250
rect 494 259 501 261
rect 494 257 496 259
rect 498 257 501 259
rect 494 252 501 257
rect 494 250 496 252
rect 498 250 501 252
rect 494 248 501 250
rect 483 243 486 245
rect 488 243 490 245
rect 483 241 490 243
rect 496 241 501 248
rect 503 260 509 269
rect 555 260 561 269
rect 503 252 511 260
rect 503 250 506 252
rect 508 250 511 252
rect 503 245 511 250
rect 503 243 506 245
rect 508 243 511 245
rect 503 241 511 243
rect 513 258 521 260
rect 513 256 516 258
rect 518 256 521 258
rect 513 251 521 256
rect 513 249 516 251
rect 518 249 521 251
rect 513 241 521 249
rect 523 252 530 260
rect 523 250 526 252
rect 528 250 530 252
rect 523 245 530 250
rect 523 243 526 245
rect 528 243 530 245
rect 523 241 530 243
rect 534 252 541 260
rect 534 250 536 252
rect 538 250 541 252
rect 534 245 541 250
rect 534 243 536 245
rect 538 243 541 245
rect 534 241 541 243
rect 543 258 551 260
rect 543 256 546 258
rect 548 256 551 258
rect 543 251 551 256
rect 543 249 546 251
rect 548 249 551 251
rect 543 241 551 249
rect 553 252 561 260
rect 553 250 556 252
rect 558 250 561 252
rect 553 245 561 250
rect 553 243 556 245
rect 558 243 561 245
rect 553 241 561 243
rect 563 261 568 269
rect 563 259 570 261
rect 595 260 601 269
rect 563 257 566 259
rect 568 257 570 259
rect 563 252 570 257
rect 563 250 566 252
rect 568 250 570 252
rect 563 248 570 250
rect 574 252 581 260
rect 574 250 576 252
rect 578 250 581 252
rect 563 241 568 248
rect 574 245 581 250
rect 574 243 576 245
rect 578 243 581 245
rect 574 241 581 243
rect 583 258 591 260
rect 583 256 586 258
rect 588 256 591 258
rect 583 251 591 256
rect 583 249 586 251
rect 588 249 591 251
rect 583 241 591 249
rect 593 252 601 260
rect 593 250 596 252
rect 598 250 601 252
rect 593 245 601 250
rect 593 243 596 245
rect 598 243 601 245
rect 593 241 601 243
rect 603 261 608 269
rect 615 267 622 269
rect 615 265 617 267
rect 619 265 622 267
rect 603 259 610 261
rect 603 257 606 259
rect 608 257 610 259
rect 603 252 610 257
rect 615 260 622 265
rect 615 258 617 260
rect 619 258 622 260
rect 615 256 622 258
rect 603 250 606 252
rect 608 250 610 252
rect 603 248 610 250
rect 603 241 608 248
rect 617 241 622 256
rect 624 252 632 269
rect 624 250 627 252
rect 629 250 632 252
rect 624 245 632 250
rect 624 243 627 245
rect 629 243 632 245
rect 624 241 632 243
rect 634 260 642 269
rect 634 258 637 260
rect 639 258 642 260
rect 634 253 642 258
rect 634 251 637 253
rect 639 251 642 253
rect 634 241 642 251
rect 644 252 660 269
rect 644 250 649 252
rect 651 250 660 252
rect 644 245 660 250
rect 644 243 649 245
rect 651 244 660 245
rect 662 244 667 269
rect 669 266 674 269
rect 669 264 677 266
rect 669 262 672 264
rect 674 262 677 264
rect 669 253 677 262
rect 679 253 690 266
rect 669 244 674 253
rect 681 245 690 253
rect 651 243 658 244
rect 644 241 658 243
rect 681 243 684 245
rect 686 243 690 245
rect 681 241 690 243
rect 692 264 699 266
rect 692 262 695 264
rect 697 262 699 264
rect 692 257 699 262
rect 692 255 695 257
rect 697 255 699 257
rect 692 253 699 255
rect 692 241 697 253
rect 29 230 36 232
rect 29 229 31 230
rect 20 223 25 229
rect 18 221 25 223
rect 18 219 20 221
rect 22 219 25 221
rect 18 214 25 219
rect 18 212 20 214
rect 22 212 25 214
rect 18 210 25 212
rect 20 201 25 210
rect 27 228 31 229
rect 33 229 36 230
rect 33 228 38 229
rect 27 201 38 228
rect 40 201 45 229
rect 47 223 52 229
rect 47 221 54 223
rect 47 219 50 221
rect 52 219 54 221
rect 47 217 54 219
rect 47 201 52 217
rect 61 214 66 229
rect 59 212 66 214
rect 59 210 61 212
rect 63 210 66 212
rect 59 205 66 210
rect 59 203 61 205
rect 63 203 66 205
rect 59 201 66 203
rect 68 227 76 229
rect 68 225 71 227
rect 73 225 76 227
rect 68 220 76 225
rect 68 218 71 220
rect 73 218 76 220
rect 68 201 76 218
rect 78 219 86 229
rect 78 217 81 219
rect 83 217 86 219
rect 78 212 86 217
rect 78 210 81 212
rect 83 210 86 212
rect 78 201 86 210
rect 88 227 102 229
rect 88 225 93 227
rect 95 226 102 227
rect 125 227 134 229
rect 95 225 104 226
rect 88 220 104 225
rect 88 218 93 220
rect 95 218 104 220
rect 88 201 104 218
rect 106 201 111 226
rect 113 217 118 226
rect 125 225 128 227
rect 130 225 134 227
rect 125 217 134 225
rect 113 208 121 217
rect 113 206 116 208
rect 118 206 121 208
rect 113 204 121 206
rect 123 204 134 217
rect 136 217 141 229
rect 136 215 143 217
rect 136 213 139 215
rect 141 213 143 215
rect 162 214 167 229
rect 136 208 143 213
rect 136 206 139 208
rect 141 206 143 208
rect 136 204 143 206
rect 160 212 167 214
rect 160 210 162 212
rect 164 210 167 212
rect 160 205 167 210
rect 113 201 118 204
rect 160 203 162 205
rect 164 203 167 205
rect 160 201 167 203
rect 169 227 177 229
rect 169 225 172 227
rect 174 225 177 227
rect 169 220 177 225
rect 169 218 172 220
rect 174 218 177 220
rect 169 201 177 218
rect 179 219 187 229
rect 179 217 182 219
rect 184 217 187 219
rect 179 212 187 217
rect 179 210 182 212
rect 184 210 187 212
rect 179 201 187 210
rect 189 227 203 229
rect 189 225 194 227
rect 196 226 203 227
rect 226 227 235 229
rect 196 225 205 226
rect 189 220 205 225
rect 189 218 194 220
rect 196 218 205 220
rect 189 201 205 218
rect 207 201 212 226
rect 214 217 219 226
rect 226 225 229 227
rect 231 225 235 227
rect 226 217 235 225
rect 214 208 222 217
rect 214 206 217 208
rect 219 206 222 208
rect 214 204 222 206
rect 224 204 235 217
rect 237 217 242 229
rect 237 215 244 217
rect 237 213 240 215
rect 242 213 244 215
rect 264 214 269 229
rect 237 208 244 213
rect 237 206 240 208
rect 242 206 244 208
rect 237 204 244 206
rect 262 212 269 214
rect 262 210 264 212
rect 266 210 269 212
rect 262 205 269 210
rect 214 201 219 204
rect 262 203 264 205
rect 266 203 269 205
rect 262 201 269 203
rect 271 227 279 229
rect 271 225 274 227
rect 276 225 279 227
rect 271 220 279 225
rect 271 218 274 220
rect 276 218 279 220
rect 271 201 279 218
rect 281 219 289 229
rect 281 217 284 219
rect 286 217 289 219
rect 281 212 289 217
rect 281 210 284 212
rect 286 210 289 212
rect 281 201 289 210
rect 291 227 305 229
rect 291 225 296 227
rect 298 226 305 227
rect 373 230 380 232
rect 373 229 375 230
rect 328 227 337 229
rect 298 225 307 226
rect 291 220 307 225
rect 291 218 296 220
rect 298 218 307 220
rect 291 201 307 218
rect 309 201 314 226
rect 316 217 321 226
rect 328 225 331 227
rect 333 225 337 227
rect 328 217 337 225
rect 316 208 324 217
rect 316 206 319 208
rect 321 206 324 208
rect 316 204 324 206
rect 326 204 337 217
rect 339 217 344 229
rect 364 223 369 229
rect 362 221 369 223
rect 362 219 364 221
rect 366 219 369 221
rect 339 215 346 217
rect 339 213 342 215
rect 344 213 346 215
rect 339 208 346 213
rect 362 214 369 219
rect 362 212 364 214
rect 366 212 369 214
rect 362 210 369 212
rect 339 206 342 208
rect 344 206 346 208
rect 339 204 346 206
rect 316 201 321 204
rect 364 201 369 210
rect 371 228 375 229
rect 377 229 380 230
rect 377 228 382 229
rect 371 201 382 228
rect 384 201 389 229
rect 391 223 396 229
rect 391 221 398 223
rect 391 219 394 221
rect 396 219 398 221
rect 391 217 398 219
rect 391 201 396 217
rect 417 214 422 229
rect 415 212 422 214
rect 415 210 417 212
rect 419 210 422 212
rect 415 205 422 210
rect 415 203 417 205
rect 419 203 422 205
rect 415 201 422 203
rect 424 227 432 229
rect 424 225 427 227
rect 429 225 432 227
rect 424 220 432 225
rect 424 218 427 220
rect 429 218 432 220
rect 424 201 432 218
rect 434 219 442 229
rect 434 217 437 219
rect 439 217 442 219
rect 434 212 442 217
rect 434 210 437 212
rect 439 210 442 212
rect 434 201 442 210
rect 444 227 458 229
rect 444 225 449 227
rect 451 226 458 227
rect 481 227 490 229
rect 451 225 460 226
rect 444 220 460 225
rect 444 218 449 220
rect 451 218 460 220
rect 444 201 460 218
rect 462 201 467 226
rect 469 217 474 226
rect 481 225 484 227
rect 486 225 490 227
rect 481 217 490 225
rect 469 208 477 217
rect 469 206 472 208
rect 474 206 477 208
rect 469 204 477 206
rect 479 204 490 217
rect 492 217 497 229
rect 492 215 499 217
rect 492 213 495 215
rect 497 213 499 215
rect 518 214 523 229
rect 492 208 499 213
rect 492 206 495 208
rect 497 206 499 208
rect 492 204 499 206
rect 516 212 523 214
rect 516 210 518 212
rect 520 210 523 212
rect 516 205 523 210
rect 469 201 474 204
rect 516 203 518 205
rect 520 203 523 205
rect 516 201 523 203
rect 525 227 533 229
rect 525 225 528 227
rect 530 225 533 227
rect 525 220 533 225
rect 525 218 528 220
rect 530 218 533 220
rect 525 201 533 218
rect 535 219 543 229
rect 535 217 538 219
rect 540 217 543 219
rect 535 212 543 217
rect 535 210 538 212
rect 540 210 543 212
rect 535 201 543 210
rect 545 227 559 229
rect 545 225 550 227
rect 552 226 559 227
rect 582 227 591 229
rect 552 225 561 226
rect 545 220 561 225
rect 545 218 550 220
rect 552 218 561 220
rect 545 201 561 218
rect 563 201 568 226
rect 570 217 575 226
rect 582 225 585 227
rect 587 225 591 227
rect 582 217 591 225
rect 570 208 578 217
rect 570 206 573 208
rect 575 206 578 208
rect 570 204 578 206
rect 580 204 591 217
rect 593 217 598 229
rect 593 215 600 217
rect 593 213 596 215
rect 598 213 600 215
rect 617 214 622 229
rect 593 208 600 213
rect 593 206 596 208
rect 598 206 600 208
rect 593 204 600 206
rect 615 212 622 214
rect 615 210 617 212
rect 619 210 622 212
rect 615 205 622 210
rect 570 201 575 204
rect 615 203 617 205
rect 619 203 622 205
rect 615 201 622 203
rect 624 227 632 229
rect 624 225 627 227
rect 629 225 632 227
rect 624 220 632 225
rect 624 218 627 220
rect 629 218 632 220
rect 624 201 632 218
rect 634 219 642 229
rect 634 217 637 219
rect 639 217 642 219
rect 634 212 642 217
rect 634 210 637 212
rect 639 210 642 212
rect 634 201 642 210
rect 644 227 658 229
rect 644 225 649 227
rect 651 226 658 227
rect 681 227 690 229
rect 651 225 660 226
rect 644 220 660 225
rect 644 218 649 220
rect 651 218 660 220
rect 644 201 660 218
rect 662 201 667 226
rect 669 217 674 226
rect 681 225 684 227
rect 686 225 690 227
rect 681 217 690 225
rect 669 208 677 217
rect 669 206 672 208
rect 674 206 677 208
rect 669 204 677 206
rect 679 204 690 217
rect 692 217 697 229
rect 692 215 699 217
rect 692 213 695 215
rect 697 213 699 215
rect 692 208 699 213
rect 692 206 695 208
rect 697 206 699 208
rect 692 204 699 206
rect 669 201 674 204
rect 20 123 27 125
rect 20 121 22 123
rect 24 121 27 123
rect 20 116 27 121
rect 20 114 22 116
rect 24 114 27 116
rect 20 112 27 114
rect 22 97 27 112
rect 29 108 37 125
rect 29 106 32 108
rect 34 106 37 108
rect 29 101 37 106
rect 29 99 32 101
rect 34 99 37 101
rect 29 97 37 99
rect 39 116 47 125
rect 39 114 42 116
rect 44 114 47 116
rect 39 109 47 114
rect 39 107 42 109
rect 44 107 47 109
rect 39 97 47 107
rect 49 108 65 125
rect 49 106 54 108
rect 56 106 65 108
rect 49 101 65 106
rect 49 99 54 101
rect 56 100 65 101
rect 67 100 72 125
rect 74 122 79 125
rect 74 120 82 122
rect 74 118 77 120
rect 79 118 82 120
rect 74 109 82 118
rect 84 109 95 122
rect 74 100 79 109
rect 86 101 95 109
rect 56 99 63 100
rect 49 97 63 99
rect 86 99 89 101
rect 91 99 95 101
rect 86 97 95 99
rect 97 120 104 122
rect 97 118 100 120
rect 102 118 104 120
rect 97 113 104 118
rect 110 116 115 125
rect 97 111 100 113
rect 102 111 104 113
rect 97 109 104 111
rect 108 114 115 116
rect 108 112 110 114
rect 112 112 115 114
rect 97 97 102 109
rect 108 107 115 112
rect 108 105 110 107
rect 112 105 115 107
rect 108 103 115 105
rect 110 97 115 103
rect 117 98 128 125
rect 117 97 121 98
rect 119 96 121 97
rect 123 97 128 98
rect 130 97 135 125
rect 137 109 142 125
rect 161 123 168 125
rect 161 121 163 123
rect 165 121 168 123
rect 161 116 168 121
rect 161 114 163 116
rect 165 114 168 116
rect 161 112 168 114
rect 137 107 144 109
rect 137 105 140 107
rect 142 105 144 107
rect 137 103 144 105
rect 137 97 142 103
rect 163 97 168 112
rect 170 108 178 125
rect 170 106 173 108
rect 175 106 178 108
rect 170 101 178 106
rect 170 99 173 101
rect 175 99 178 101
rect 170 97 178 99
rect 180 116 188 125
rect 180 114 183 116
rect 185 114 188 116
rect 180 109 188 114
rect 180 107 183 109
rect 185 107 188 109
rect 180 97 188 107
rect 190 108 206 125
rect 190 106 195 108
rect 197 106 206 108
rect 190 101 206 106
rect 190 99 195 101
rect 197 100 206 101
rect 208 100 213 125
rect 215 122 220 125
rect 286 122 291 125
rect 215 120 223 122
rect 215 118 218 120
rect 220 118 223 120
rect 215 109 223 118
rect 225 109 236 122
rect 215 100 220 109
rect 227 101 236 109
rect 197 99 204 100
rect 190 97 204 99
rect 123 96 126 97
rect 119 94 126 96
rect 227 99 230 101
rect 232 99 236 101
rect 227 97 236 99
rect 238 120 245 122
rect 238 118 241 120
rect 243 118 245 120
rect 238 113 245 118
rect 238 111 241 113
rect 243 111 245 113
rect 238 109 245 111
rect 261 120 268 122
rect 261 118 263 120
rect 265 118 268 120
rect 261 113 268 118
rect 261 111 263 113
rect 265 111 268 113
rect 261 109 268 111
rect 238 97 243 109
rect 263 97 268 109
rect 270 109 281 122
rect 283 120 291 122
rect 283 118 286 120
rect 288 118 291 120
rect 283 109 291 118
rect 270 101 279 109
rect 270 99 274 101
rect 276 99 279 101
rect 286 100 291 109
rect 293 100 298 125
rect 300 108 316 125
rect 300 106 309 108
rect 311 106 316 108
rect 300 101 316 106
rect 300 100 309 101
rect 270 97 279 99
rect 302 99 309 100
rect 311 99 316 101
rect 302 97 316 99
rect 318 116 326 125
rect 318 114 321 116
rect 323 114 326 116
rect 318 109 326 114
rect 318 107 321 109
rect 323 107 326 109
rect 318 97 326 107
rect 328 108 336 125
rect 328 106 331 108
rect 333 106 336 108
rect 328 101 336 106
rect 328 99 331 101
rect 333 99 336 101
rect 328 97 336 99
rect 338 123 345 125
rect 338 121 341 123
rect 343 121 345 123
rect 338 116 345 121
rect 364 116 369 125
rect 338 114 341 116
rect 343 114 345 116
rect 338 112 345 114
rect 362 114 369 116
rect 362 112 364 114
rect 366 112 369 114
rect 338 97 343 112
rect 362 107 369 112
rect 362 105 364 107
rect 366 105 369 107
rect 362 103 369 105
rect 364 97 369 103
rect 371 98 382 125
rect 371 97 375 98
rect 373 96 375 97
rect 377 97 382 98
rect 384 97 389 125
rect 391 109 396 125
rect 415 123 422 125
rect 415 121 417 123
rect 419 121 422 123
rect 415 116 422 121
rect 415 114 417 116
rect 419 114 422 116
rect 415 112 422 114
rect 391 107 398 109
rect 391 105 394 107
rect 396 105 398 107
rect 391 103 398 105
rect 391 97 396 103
rect 417 97 422 112
rect 424 108 432 125
rect 424 106 427 108
rect 429 106 432 108
rect 424 101 432 106
rect 424 99 427 101
rect 429 99 432 101
rect 424 97 432 99
rect 434 116 442 125
rect 434 114 437 116
rect 439 114 442 116
rect 434 109 442 114
rect 434 107 437 109
rect 439 107 442 109
rect 434 97 442 107
rect 444 108 460 125
rect 444 106 449 108
rect 451 106 460 108
rect 444 101 460 106
rect 444 99 449 101
rect 451 100 460 101
rect 462 100 467 125
rect 469 122 474 125
rect 516 123 523 125
rect 469 120 477 122
rect 469 118 472 120
rect 474 118 477 120
rect 469 109 477 118
rect 479 109 490 122
rect 469 100 474 109
rect 481 101 490 109
rect 451 99 458 100
rect 444 97 458 99
rect 377 96 380 97
rect 373 94 380 96
rect 481 99 484 101
rect 486 99 490 101
rect 481 97 490 99
rect 492 120 499 122
rect 492 118 495 120
rect 497 118 499 120
rect 492 113 499 118
rect 492 111 495 113
rect 497 111 499 113
rect 516 121 518 123
rect 520 121 523 123
rect 516 116 523 121
rect 516 114 518 116
rect 520 114 523 116
rect 516 112 523 114
rect 492 109 499 111
rect 492 97 497 109
rect 518 97 523 112
rect 525 108 533 125
rect 525 106 528 108
rect 530 106 533 108
rect 525 101 533 106
rect 525 99 528 101
rect 530 99 533 101
rect 525 97 533 99
rect 535 116 543 125
rect 535 114 538 116
rect 540 114 543 116
rect 535 109 543 114
rect 535 107 538 109
rect 540 107 543 109
rect 535 97 543 107
rect 545 108 561 125
rect 545 106 550 108
rect 552 106 561 108
rect 545 101 561 106
rect 545 99 550 101
rect 552 100 561 101
rect 563 100 568 125
rect 570 122 575 125
rect 615 123 622 125
rect 570 120 578 122
rect 570 118 573 120
rect 575 118 578 120
rect 570 109 578 118
rect 580 109 591 122
rect 570 100 575 109
rect 582 101 591 109
rect 552 99 559 100
rect 545 97 559 99
rect 582 99 585 101
rect 587 99 591 101
rect 582 97 591 99
rect 593 120 600 122
rect 593 118 596 120
rect 598 118 600 120
rect 593 113 600 118
rect 593 111 596 113
rect 598 111 600 113
rect 615 121 617 123
rect 619 121 622 123
rect 615 116 622 121
rect 615 114 617 116
rect 619 114 622 116
rect 615 112 622 114
rect 593 109 600 111
rect 593 97 598 109
rect 617 97 622 112
rect 624 108 632 125
rect 624 106 627 108
rect 629 106 632 108
rect 624 101 632 106
rect 624 99 627 101
rect 629 99 632 101
rect 624 97 632 99
rect 634 116 642 125
rect 634 114 637 116
rect 639 114 642 116
rect 634 109 642 114
rect 634 107 637 109
rect 639 107 642 109
rect 634 97 642 107
rect 644 108 660 125
rect 644 106 649 108
rect 651 106 660 108
rect 644 101 660 106
rect 644 99 649 101
rect 651 100 660 101
rect 662 100 667 125
rect 669 122 674 125
rect 669 120 677 122
rect 669 118 672 120
rect 674 118 677 120
rect 669 109 677 118
rect 679 109 690 122
rect 669 100 674 109
rect 681 101 690 109
rect 651 99 658 100
rect 644 97 658 99
rect 681 99 684 101
rect 686 99 690 101
rect 681 97 690 99
rect 692 120 699 122
rect 692 118 695 120
rect 697 118 699 120
rect 692 113 699 118
rect 692 111 695 113
rect 697 111 699 113
rect 692 109 699 111
rect 692 97 697 109
rect 29 86 36 88
rect 29 85 31 86
rect 20 79 25 85
rect 18 77 25 79
rect 18 75 20 77
rect 22 75 25 77
rect 18 70 25 75
rect 18 68 20 70
rect 22 68 25 70
rect 18 66 25 68
rect 20 57 25 66
rect 27 84 31 85
rect 33 85 36 86
rect 33 84 38 85
rect 27 57 38 84
rect 40 57 45 85
rect 47 79 52 85
rect 47 77 54 79
rect 47 75 50 77
rect 52 75 54 77
rect 47 73 54 75
rect 47 57 52 73
rect 61 70 66 85
rect 59 68 66 70
rect 59 66 61 68
rect 63 66 66 68
rect 59 61 66 66
rect 59 59 61 61
rect 63 59 66 61
rect 59 57 66 59
rect 68 83 76 85
rect 68 81 71 83
rect 73 81 76 83
rect 68 76 76 81
rect 68 74 71 76
rect 73 74 76 76
rect 68 57 76 74
rect 78 75 86 85
rect 78 73 81 75
rect 83 73 86 75
rect 78 68 86 73
rect 78 66 81 68
rect 83 66 86 68
rect 78 57 86 66
rect 88 83 102 85
rect 88 81 93 83
rect 95 82 102 83
rect 125 83 134 85
rect 95 81 104 82
rect 88 76 104 81
rect 88 74 93 76
rect 95 74 104 76
rect 88 57 104 74
rect 106 57 111 82
rect 113 73 118 82
rect 125 81 128 83
rect 130 81 134 83
rect 125 73 134 81
rect 113 64 121 73
rect 113 62 116 64
rect 118 62 121 64
rect 113 60 121 62
rect 123 60 134 73
rect 136 73 141 85
rect 136 71 143 73
rect 136 69 139 71
rect 141 69 143 71
rect 162 70 167 85
rect 136 64 143 69
rect 136 62 139 64
rect 141 62 143 64
rect 136 60 143 62
rect 160 68 167 70
rect 160 66 162 68
rect 164 66 167 68
rect 160 61 167 66
rect 113 57 118 60
rect 160 59 162 61
rect 164 59 167 61
rect 160 57 167 59
rect 169 83 177 85
rect 169 81 172 83
rect 174 81 177 83
rect 169 76 177 81
rect 169 74 172 76
rect 174 74 177 76
rect 169 57 177 74
rect 179 75 187 85
rect 179 73 182 75
rect 184 73 187 75
rect 179 68 187 73
rect 179 66 182 68
rect 184 66 187 68
rect 179 57 187 66
rect 189 83 203 85
rect 189 81 194 83
rect 196 82 203 83
rect 226 83 235 85
rect 196 81 205 82
rect 189 76 205 81
rect 189 74 194 76
rect 196 74 205 76
rect 189 57 205 74
rect 207 57 212 82
rect 214 73 219 82
rect 226 81 229 83
rect 231 81 235 83
rect 226 73 235 81
rect 214 64 222 73
rect 214 62 217 64
rect 219 62 222 64
rect 214 60 222 62
rect 224 60 235 73
rect 237 73 242 85
rect 237 71 244 73
rect 237 69 240 71
rect 242 69 244 71
rect 263 70 268 85
rect 237 64 244 69
rect 237 62 240 64
rect 242 62 244 64
rect 237 60 244 62
rect 261 68 268 70
rect 261 66 263 68
rect 265 66 268 68
rect 261 61 268 66
rect 214 57 219 60
rect 261 59 263 61
rect 265 59 268 61
rect 261 57 268 59
rect 270 83 278 85
rect 270 81 273 83
rect 275 81 278 83
rect 270 76 278 81
rect 270 74 273 76
rect 275 74 278 76
rect 270 57 278 74
rect 280 75 288 85
rect 280 73 283 75
rect 285 73 288 75
rect 280 68 288 73
rect 280 66 283 68
rect 285 66 288 68
rect 280 57 288 66
rect 290 83 304 85
rect 290 81 295 83
rect 297 82 304 83
rect 372 86 379 88
rect 372 85 374 86
rect 327 83 336 85
rect 297 81 306 82
rect 290 76 306 81
rect 290 74 295 76
rect 297 74 306 76
rect 290 57 306 74
rect 308 57 313 82
rect 315 73 320 82
rect 327 81 330 83
rect 332 81 336 83
rect 327 73 336 81
rect 315 64 323 73
rect 315 62 318 64
rect 320 62 323 64
rect 315 60 323 62
rect 325 60 336 73
rect 338 73 343 85
rect 363 79 368 85
rect 361 77 368 79
rect 361 75 363 77
rect 365 75 368 77
rect 338 71 345 73
rect 338 69 341 71
rect 343 69 345 71
rect 338 64 345 69
rect 361 70 368 75
rect 361 68 363 70
rect 365 68 368 70
rect 361 66 368 68
rect 338 62 341 64
rect 343 62 345 64
rect 338 60 345 62
rect 315 57 320 60
rect 363 57 368 66
rect 370 84 374 85
rect 376 85 379 86
rect 376 84 381 85
rect 370 57 381 84
rect 383 57 388 85
rect 390 79 395 85
rect 390 77 397 79
rect 390 75 393 77
rect 395 75 397 77
rect 390 73 397 75
rect 390 57 395 73
rect 416 70 421 85
rect 414 68 421 70
rect 414 66 416 68
rect 418 66 421 68
rect 414 61 421 66
rect 414 59 416 61
rect 418 59 421 61
rect 414 57 421 59
rect 423 83 431 85
rect 423 81 426 83
rect 428 81 431 83
rect 423 76 431 81
rect 423 74 426 76
rect 428 74 431 76
rect 423 57 431 74
rect 433 75 441 85
rect 433 73 436 75
rect 438 73 441 75
rect 433 68 441 73
rect 433 66 436 68
rect 438 66 441 68
rect 433 57 441 66
rect 443 83 457 85
rect 443 81 448 83
rect 450 82 457 83
rect 480 83 489 85
rect 450 81 459 82
rect 443 76 459 81
rect 443 74 448 76
rect 450 74 459 76
rect 443 57 459 74
rect 461 57 466 82
rect 468 73 473 82
rect 480 81 483 83
rect 485 81 489 83
rect 480 73 489 81
rect 468 64 476 73
rect 468 62 471 64
rect 473 62 476 64
rect 468 60 476 62
rect 478 60 489 73
rect 491 73 496 85
rect 491 71 498 73
rect 491 69 494 71
rect 496 69 498 71
rect 517 70 522 85
rect 491 64 498 69
rect 491 62 494 64
rect 496 62 498 64
rect 491 60 498 62
rect 515 68 522 70
rect 515 66 517 68
rect 519 66 522 68
rect 515 61 522 66
rect 468 57 473 60
rect 515 59 517 61
rect 519 59 522 61
rect 515 57 522 59
rect 524 83 532 85
rect 524 81 527 83
rect 529 81 532 83
rect 524 76 532 81
rect 524 74 527 76
rect 529 74 532 76
rect 524 57 532 74
rect 534 75 542 85
rect 534 73 537 75
rect 539 73 542 75
rect 534 68 542 73
rect 534 66 537 68
rect 539 66 542 68
rect 534 57 542 66
rect 544 83 558 85
rect 544 81 549 83
rect 551 82 558 83
rect 581 83 590 85
rect 551 81 560 82
rect 544 76 560 81
rect 544 74 549 76
rect 551 74 560 76
rect 544 57 560 74
rect 562 57 567 82
rect 569 73 574 82
rect 581 81 584 83
rect 586 81 590 83
rect 581 73 590 81
rect 569 64 577 73
rect 569 62 572 64
rect 574 62 577 64
rect 569 60 577 62
rect 579 60 590 73
rect 592 73 597 85
rect 592 71 599 73
rect 592 69 595 71
rect 597 69 599 71
rect 616 70 621 85
rect 592 64 599 69
rect 592 62 595 64
rect 597 62 599 64
rect 592 60 599 62
rect 614 68 621 70
rect 614 66 616 68
rect 618 66 621 68
rect 614 61 621 66
rect 569 57 574 60
rect 614 59 616 61
rect 618 59 621 61
rect 614 57 621 59
rect 623 83 631 85
rect 623 81 626 83
rect 628 81 631 83
rect 623 76 631 81
rect 623 74 626 76
rect 628 74 631 76
rect 623 57 631 74
rect 633 75 641 85
rect 633 73 636 75
rect 638 73 641 75
rect 633 68 641 73
rect 633 66 636 68
rect 638 66 641 68
rect 633 57 641 66
rect 643 83 657 85
rect 643 81 648 83
rect 650 82 657 83
rect 680 83 689 85
rect 650 81 659 82
rect 643 76 659 81
rect 643 74 648 76
rect 650 74 659 76
rect 643 57 659 74
rect 661 57 666 82
rect 668 73 673 82
rect 680 81 683 83
rect 685 81 689 83
rect 680 73 689 81
rect 668 64 676 73
rect 668 62 671 64
rect 673 62 676 64
rect 668 60 676 62
rect 678 60 689 73
rect 691 73 696 85
rect 691 71 698 73
rect 691 69 694 71
rect 696 69 698 71
rect 691 64 698 69
rect 691 62 694 64
rect 696 62 698 64
rect 691 60 698 62
rect 668 57 673 60
<< alu1 >>
rect 14 375 703 379
rect -1 371 703 375
rect -1 243 3 371
rect 49 364 54 366
rect 49 362 50 364
rect 52 362 54 364
rect 18 349 22 358
rect 49 357 54 362
rect 89 364 94 366
rect 89 362 90 364
rect 92 362 94 364
rect 49 355 50 357
rect 52 355 54 357
rect 49 353 54 355
rect 18 348 31 349
rect 18 346 23 348
rect 25 346 28 348
rect 30 346 31 348
rect 18 345 31 346
rect 25 340 39 341
rect 25 338 33 340
rect 35 338 39 340
rect 25 337 39 338
rect 25 331 30 337
rect 25 329 26 331
rect 28 329 30 331
rect 25 328 30 329
rect 50 331 54 353
rect 58 349 62 358
rect 89 357 94 362
rect 170 361 183 365
rect 89 355 90 357
rect 92 355 94 357
rect 89 353 94 355
rect 58 348 71 349
rect 58 346 59 348
rect 61 346 63 348
rect 65 346 71 348
rect 58 345 71 346
rect 52 329 54 331
rect 50 326 54 329
rect 65 340 79 341
rect 65 338 73 340
rect 75 338 79 340
rect 65 337 79 338
rect 65 331 70 337
rect 65 329 66 331
rect 68 329 70 331
rect 65 328 70 329
rect 42 323 54 326
rect 90 331 94 353
rect 92 329 94 331
rect 90 326 94 329
rect 42 321 50 323
rect 52 321 54 323
rect 82 323 94 326
rect 82 321 90 323
rect 92 321 94 323
rect 98 356 104 358
rect 178 359 183 361
rect 178 357 179 359
rect 181 357 183 359
rect 98 354 101 356
rect 103 354 104 356
rect 98 349 104 354
rect 98 347 101 349
rect 103 347 104 349
rect 98 345 104 347
rect 98 325 102 345
rect 114 348 152 349
rect 114 346 115 348
rect 117 346 152 348
rect 114 345 152 346
rect 147 342 152 345
rect 122 340 137 341
rect 122 338 126 340
rect 128 338 133 340
rect 135 338 137 340
rect 122 337 137 338
rect 147 340 155 342
rect 147 338 152 340
rect 154 338 155 340
rect 131 331 135 337
rect 147 336 155 338
rect 178 352 183 357
rect 178 350 179 352
rect 181 350 183 352
rect 178 348 183 350
rect 131 329 132 331
rect 134 329 135 331
rect 131 328 135 329
rect 98 324 120 325
rect 98 322 101 324
rect 103 322 117 324
rect 119 322 120 324
rect 98 321 120 322
rect 179 326 183 348
rect 178 324 183 326
rect 178 322 179 324
rect 181 322 183 324
rect 42 320 54 321
rect 82 320 94 321
rect 178 320 183 322
rect 195 361 208 365
rect 284 364 289 366
rect 284 362 286 364
rect 288 362 289 364
rect 195 359 200 361
rect 195 357 197 359
rect 199 357 200 359
rect 195 352 200 357
rect 195 350 197 352
rect 199 350 200 352
rect 195 348 200 350
rect 195 326 199 348
rect 226 348 264 349
rect 226 346 261 348
rect 263 346 264 348
rect 226 345 264 346
rect 226 342 231 345
rect 223 340 231 342
rect 223 338 224 340
rect 226 338 231 340
rect 223 336 231 338
rect 241 340 256 341
rect 241 338 243 340
rect 245 338 250 340
rect 252 338 256 340
rect 241 337 256 338
rect 195 324 200 326
rect 243 331 247 337
rect 274 356 280 358
rect 274 354 275 356
rect 277 354 280 356
rect 274 349 280 354
rect 274 347 275 349
rect 277 347 280 349
rect 274 345 280 347
rect 243 329 244 331
rect 246 329 247 331
rect 243 328 247 329
rect 276 325 280 345
rect 195 322 197 324
rect 199 322 200 324
rect 195 320 200 322
rect 258 324 280 325
rect 258 322 259 324
rect 261 322 275 324
rect 277 322 280 324
rect 258 321 280 322
rect 284 357 289 362
rect 324 364 329 366
rect 324 362 326 364
rect 328 362 329 364
rect 284 355 286 357
rect 288 355 289 357
rect 284 353 289 355
rect 284 331 288 353
rect 316 349 320 358
rect 307 348 320 349
rect 307 346 313 348
rect 315 346 317 348
rect 319 346 320 348
rect 307 345 320 346
rect 324 357 329 362
rect 365 361 378 365
rect 454 364 459 366
rect 454 362 456 364
rect 458 362 459 364
rect 365 359 370 361
rect 324 355 326 357
rect 328 355 329 357
rect 324 353 329 355
rect 299 340 313 341
rect 299 338 303 340
rect 305 338 313 340
rect 299 337 313 338
rect 284 329 286 331
rect 284 326 288 329
rect 284 323 296 326
rect 284 321 286 323
rect 288 321 296 323
rect 308 331 313 337
rect 308 329 310 331
rect 312 329 313 331
rect 308 328 313 329
rect 324 331 328 353
rect 356 349 360 358
rect 347 348 360 349
rect 347 346 348 348
rect 350 346 353 348
rect 355 346 360 348
rect 347 345 360 346
rect 365 357 367 359
rect 369 357 370 359
rect 365 352 370 357
rect 365 350 367 352
rect 369 350 370 352
rect 365 348 370 350
rect 339 340 353 341
rect 339 338 343 340
rect 345 338 353 340
rect 339 337 353 338
rect 324 329 326 331
rect 324 326 328 329
rect 324 323 336 326
rect 324 321 326 323
rect 328 321 336 323
rect 348 331 353 337
rect 348 329 350 331
rect 352 329 353 331
rect 348 328 353 329
rect 365 326 369 348
rect 396 348 434 349
rect 396 346 431 348
rect 433 346 434 348
rect 396 345 434 346
rect 396 342 401 345
rect 393 340 401 342
rect 393 338 394 340
rect 396 338 401 340
rect 393 336 401 338
rect 411 340 426 341
rect 411 338 413 340
rect 415 338 420 340
rect 422 338 426 340
rect 411 337 426 338
rect 365 324 370 326
rect 413 331 417 337
rect 444 356 450 358
rect 444 354 445 356
rect 447 354 450 356
rect 444 349 450 354
rect 444 347 445 349
rect 447 347 450 349
rect 444 345 450 347
rect 413 329 414 331
rect 416 329 417 331
rect 413 328 417 329
rect 446 325 450 345
rect 365 322 367 324
rect 369 322 370 324
rect 284 320 296 321
rect 324 320 336 321
rect 365 320 370 322
rect 428 324 450 325
rect 428 322 429 324
rect 431 322 445 324
rect 447 322 450 324
rect 428 321 450 322
rect 454 357 459 362
rect 494 364 499 366
rect 494 362 496 364
rect 498 362 499 364
rect 454 355 456 357
rect 458 355 459 357
rect 454 353 459 355
rect 454 331 458 353
rect 486 349 490 358
rect 477 348 490 349
rect 477 346 483 348
rect 485 346 487 348
rect 489 346 490 348
rect 477 345 490 346
rect 494 357 499 362
rect 565 364 570 366
rect 565 362 566 364
rect 568 362 570 364
rect 494 355 496 357
rect 498 355 499 357
rect 494 353 499 355
rect 469 340 483 341
rect 469 338 473 340
rect 475 338 483 340
rect 469 337 483 338
rect 454 329 456 331
rect 454 326 458 329
rect 454 323 466 326
rect 454 321 456 323
rect 458 321 466 323
rect 478 331 483 337
rect 478 329 480 331
rect 482 329 483 331
rect 478 328 483 329
rect 494 331 498 353
rect 526 349 530 358
rect 517 348 530 349
rect 517 346 518 348
rect 520 346 523 348
rect 525 346 530 348
rect 517 345 530 346
rect 534 349 538 358
rect 565 357 570 362
rect 605 364 610 366
rect 605 362 606 364
rect 608 362 610 364
rect 565 355 566 357
rect 568 355 570 357
rect 565 353 570 355
rect 534 348 547 349
rect 534 346 539 348
rect 541 346 544 348
rect 546 346 547 348
rect 534 345 547 346
rect 509 340 523 341
rect 509 338 513 340
rect 515 338 523 340
rect 509 337 523 338
rect 494 329 496 331
rect 494 326 498 329
rect 494 323 506 326
rect 494 321 496 323
rect 498 321 506 323
rect 518 331 523 337
rect 518 329 520 331
rect 522 329 523 331
rect 518 328 523 329
rect 541 340 555 341
rect 541 338 549 340
rect 551 338 555 340
rect 541 337 555 338
rect 541 331 546 337
rect 541 329 542 331
rect 544 329 546 331
rect 541 328 546 329
rect 566 331 570 353
rect 574 349 578 358
rect 605 357 610 362
rect 686 361 699 365
rect 605 355 606 357
rect 608 355 610 357
rect 605 353 610 355
rect 574 348 587 349
rect 574 346 575 348
rect 577 346 579 348
rect 581 346 587 348
rect 574 345 587 346
rect 568 329 570 331
rect 566 326 570 329
rect 581 340 595 341
rect 581 338 589 340
rect 591 338 595 340
rect 581 337 595 338
rect 581 331 586 337
rect 581 329 582 331
rect 584 329 586 331
rect 581 328 586 329
rect 558 323 570 326
rect 606 331 610 353
rect 608 329 610 331
rect 606 326 610 329
rect 558 321 566 323
rect 568 321 570 323
rect 598 323 610 326
rect 598 321 606 323
rect 608 321 610 323
rect 614 356 620 358
rect 694 359 699 361
rect 694 357 695 359
rect 697 357 699 359
rect 614 354 617 356
rect 619 354 620 356
rect 614 349 620 354
rect 614 347 617 349
rect 619 347 620 349
rect 614 345 620 347
rect 614 325 618 345
rect 630 348 668 349
rect 630 346 631 348
rect 633 346 668 348
rect 630 345 668 346
rect 663 342 668 345
rect 638 340 653 341
rect 638 338 642 340
rect 644 338 649 340
rect 651 338 653 340
rect 638 337 653 338
rect 663 340 671 342
rect 663 338 668 340
rect 670 338 671 340
rect 647 331 651 337
rect 663 336 671 338
rect 694 352 699 357
rect 694 350 695 352
rect 697 350 699 352
rect 694 348 699 350
rect 647 329 648 331
rect 650 329 651 331
rect 647 328 651 329
rect 614 324 636 325
rect 614 322 617 324
rect 619 322 633 324
rect 635 322 636 324
rect 614 321 636 322
rect 695 326 699 348
rect 694 324 699 326
rect 694 322 695 324
rect 697 322 699 324
rect 454 320 466 321
rect 494 320 506 321
rect 558 320 570 321
rect 598 320 610 321
rect 694 320 699 322
rect 14 314 703 315
rect 14 312 39 314
rect 41 312 79 314
rect 81 312 297 314
rect 299 312 337 314
rect 339 312 467 314
rect 469 312 507 314
rect 509 312 555 314
rect 557 312 595 314
rect 597 312 703 314
rect 14 303 703 312
rect 14 302 715 303
rect 14 300 39 302
rect 41 300 79 302
rect 81 300 297 302
rect 299 300 337 302
rect 339 300 467 302
rect 469 300 507 302
rect 509 300 555 302
rect 557 300 595 302
rect 597 300 715 302
rect 14 299 715 300
rect 42 293 54 294
rect 82 293 94 294
rect 25 285 30 286
rect 25 283 26 285
rect 28 283 30 285
rect 25 277 30 283
rect 42 291 50 293
rect 52 291 54 293
rect 42 288 54 291
rect 50 285 54 288
rect 52 283 54 285
rect 25 276 39 277
rect 25 274 33 276
rect 35 274 39 276
rect 25 273 39 274
rect 18 268 31 269
rect 18 266 23 268
rect 25 266 28 268
rect 30 266 31 268
rect 18 265 31 266
rect 50 276 54 283
rect 50 274 51 276
rect 53 274 54 276
rect 18 256 22 265
rect 50 261 54 274
rect 65 285 70 286
rect 65 283 66 285
rect 68 283 70 285
rect 65 277 70 283
rect 82 291 90 293
rect 92 291 94 293
rect 82 288 94 291
rect 90 285 94 288
rect 92 283 94 285
rect 65 276 79 277
rect 65 274 73 276
rect 75 274 79 276
rect 65 273 79 274
rect 49 259 54 261
rect 49 257 50 259
rect 52 257 54 259
rect 49 252 54 257
rect 58 268 71 269
rect 58 266 59 268
rect 61 266 63 268
rect 65 266 71 268
rect 58 265 71 266
rect 58 256 62 265
rect 90 261 94 283
rect 89 259 94 261
rect 89 257 90 259
rect 92 257 94 259
rect 49 250 50 252
rect 52 250 54 252
rect 49 248 54 250
rect 89 252 94 257
rect 98 292 120 293
rect 98 290 101 292
rect 103 290 120 292
rect 98 289 120 290
rect 178 292 183 294
rect 178 290 179 292
rect 181 290 183 292
rect 98 269 102 289
rect 98 267 104 269
rect 98 265 101 267
rect 103 265 104 267
rect 98 261 104 265
rect 98 257 100 261
rect 131 277 135 286
rect 178 288 183 290
rect 122 276 137 277
rect 122 274 123 276
rect 125 274 126 276
rect 128 274 133 276
rect 135 274 137 276
rect 122 273 137 274
rect 147 276 155 278
rect 147 274 152 276
rect 154 274 155 276
rect 147 272 155 274
rect 147 269 152 272
rect 114 268 152 269
rect 114 266 115 268
rect 117 266 152 268
rect 114 265 152 266
rect 179 266 183 288
rect 178 264 183 266
rect 178 262 179 264
rect 181 262 183 264
rect 178 257 183 262
rect 98 256 104 257
rect 178 255 179 257
rect 181 255 183 257
rect 178 253 183 255
rect 89 250 90 252
rect 92 250 94 252
rect 89 248 94 250
rect 170 249 183 253
rect 195 292 200 294
rect 284 293 296 294
rect 324 293 336 294
rect 195 290 197 292
rect 199 290 200 292
rect 195 288 200 290
rect 195 266 199 288
rect 258 292 280 293
rect 258 290 275 292
rect 277 290 280 292
rect 258 289 280 290
rect 195 264 200 266
rect 195 262 197 264
rect 199 262 200 264
rect 195 257 200 262
rect 223 276 231 278
rect 243 277 247 286
rect 223 274 224 276
rect 226 274 231 276
rect 223 272 231 274
rect 241 276 256 277
rect 241 274 243 276
rect 245 274 250 276
rect 252 274 253 276
rect 255 274 256 276
rect 241 273 256 274
rect 226 269 231 272
rect 226 268 264 269
rect 226 266 261 268
rect 263 266 264 268
rect 226 265 264 266
rect 276 269 280 289
rect 274 267 280 269
rect 274 265 275 267
rect 277 265 280 267
rect 274 260 280 265
rect 274 258 275 260
rect 277 258 280 260
rect 195 255 197 257
rect 199 255 200 257
rect 195 253 200 255
rect 274 256 280 258
rect 284 291 286 293
rect 288 291 296 293
rect 284 288 296 291
rect 324 291 326 293
rect 328 291 336 293
rect 284 285 288 288
rect 284 283 286 285
rect 284 261 288 283
rect 324 288 336 291
rect 365 292 370 294
rect 454 293 466 294
rect 494 293 506 294
rect 558 293 570 294
rect 598 293 610 294
rect 365 290 367 292
rect 369 290 370 292
rect 308 285 313 286
rect 308 283 310 285
rect 312 283 313 285
rect 308 277 313 283
rect 299 276 313 277
rect 299 274 303 276
rect 305 274 313 276
rect 299 273 313 274
rect 324 285 328 288
rect 324 283 326 285
rect 307 268 320 269
rect 307 266 313 268
rect 315 266 317 268
rect 319 266 320 268
rect 307 265 320 266
rect 284 259 289 261
rect 284 257 286 259
rect 288 257 289 259
rect 195 249 208 253
rect 284 252 289 257
rect 316 256 320 265
rect 324 261 328 283
rect 365 288 370 290
rect 348 285 353 286
rect 348 283 350 285
rect 352 283 353 285
rect 348 277 353 283
rect 339 276 353 277
rect 339 274 343 276
rect 345 274 353 276
rect 339 273 353 274
rect 347 268 360 269
rect 347 266 348 268
rect 350 266 353 268
rect 355 266 360 268
rect 347 265 360 266
rect 324 259 329 261
rect 324 257 326 259
rect 328 257 329 259
rect 284 250 286 252
rect 288 250 289 252
rect 284 248 289 250
rect 324 255 329 257
rect 324 253 326 255
rect 328 253 329 255
rect 356 256 360 265
rect 365 266 369 288
rect 428 292 450 293
rect 428 290 445 292
rect 447 290 450 292
rect 428 289 450 290
rect 365 264 370 266
rect 365 262 367 264
rect 369 262 370 264
rect 365 257 370 262
rect 393 276 401 278
rect 413 277 417 286
rect 446 284 450 289
rect 446 282 447 284
rect 449 282 450 284
rect 393 274 394 276
rect 396 274 401 276
rect 393 272 401 274
rect 411 276 426 277
rect 411 274 413 276
rect 415 274 420 276
rect 422 274 423 276
rect 425 274 426 276
rect 411 273 426 274
rect 396 269 401 272
rect 396 268 434 269
rect 396 266 431 268
rect 433 266 434 268
rect 396 265 434 266
rect 446 269 450 282
rect 444 267 450 269
rect 444 265 445 267
rect 447 265 450 267
rect 444 260 450 265
rect 444 258 445 260
rect 447 258 450 260
rect 324 252 329 253
rect 324 250 326 252
rect 328 250 329 252
rect 324 248 329 250
rect 365 255 367 257
rect 369 255 370 257
rect 365 253 370 255
rect 444 256 450 258
rect 454 291 456 293
rect 458 291 466 293
rect 454 288 466 291
rect 494 291 496 293
rect 498 291 506 293
rect 454 285 458 288
rect 454 283 456 285
rect 454 261 458 283
rect 494 288 506 291
rect 478 285 483 286
rect 478 283 480 285
rect 482 283 483 285
rect 478 277 483 283
rect 469 276 483 277
rect 469 274 473 276
rect 475 274 483 276
rect 469 273 483 274
rect 494 285 498 288
rect 494 283 496 285
rect 494 276 498 283
rect 518 285 523 286
rect 518 283 520 285
rect 522 283 523 285
rect 494 274 495 276
rect 497 274 498 276
rect 477 268 490 269
rect 477 266 483 268
rect 485 266 487 268
rect 489 266 490 268
rect 477 265 490 266
rect 454 259 459 261
rect 454 257 456 259
rect 458 257 459 259
rect 365 249 378 253
rect 454 252 459 257
rect 486 256 490 265
rect 494 261 498 274
rect 518 277 523 283
rect 509 276 523 277
rect 509 274 513 276
rect 515 274 523 276
rect 509 273 523 274
rect 541 285 546 286
rect 541 283 542 285
rect 544 283 546 285
rect 541 277 546 283
rect 558 291 566 293
rect 568 291 570 293
rect 558 288 570 291
rect 566 285 570 288
rect 568 283 570 285
rect 541 276 555 277
rect 541 274 549 276
rect 551 274 555 276
rect 541 273 555 274
rect 517 268 530 269
rect 517 266 518 268
rect 520 266 523 268
rect 525 266 530 268
rect 517 265 530 266
rect 494 259 499 261
rect 494 257 496 259
rect 498 257 499 259
rect 454 250 456 252
rect 458 250 459 252
rect 454 248 459 250
rect 494 252 499 257
rect 526 256 530 265
rect 534 268 547 269
rect 534 266 539 268
rect 541 266 544 268
rect 546 266 547 268
rect 534 265 547 266
rect 534 256 538 265
rect 566 261 570 283
rect 581 285 586 286
rect 581 283 582 285
rect 584 283 586 285
rect 581 277 586 283
rect 598 291 606 293
rect 608 291 610 293
rect 598 288 610 291
rect 606 285 610 288
rect 608 283 610 285
rect 581 276 595 277
rect 581 274 589 276
rect 591 274 595 276
rect 581 273 595 274
rect 565 259 570 261
rect 565 257 566 259
rect 568 257 570 259
rect 494 250 496 252
rect 498 250 499 252
rect 494 248 499 250
rect 565 252 570 257
rect 574 268 587 269
rect 574 266 575 268
rect 577 266 579 268
rect 581 266 587 268
rect 574 265 587 266
rect 574 256 578 265
rect 606 261 610 283
rect 605 259 610 261
rect 605 257 606 259
rect 608 257 610 259
rect 565 250 566 252
rect 568 250 570 252
rect 565 248 570 250
rect 605 252 610 257
rect 614 292 636 293
rect 614 290 617 292
rect 619 290 636 292
rect 614 289 636 290
rect 694 292 699 294
rect 694 290 695 292
rect 697 290 699 292
rect 614 269 618 289
rect 614 267 620 269
rect 614 265 617 267
rect 619 265 620 267
rect 614 260 620 265
rect 614 258 617 260
rect 619 258 620 260
rect 614 256 620 258
rect 647 277 651 286
rect 694 288 699 290
rect 638 276 653 277
rect 638 274 639 276
rect 641 274 642 276
rect 644 274 649 276
rect 651 274 653 276
rect 638 273 653 274
rect 663 276 671 278
rect 663 274 668 276
rect 670 274 671 276
rect 663 272 671 274
rect 663 269 668 272
rect 630 268 668 269
rect 630 266 631 268
rect 633 266 668 268
rect 630 265 668 266
rect 695 266 699 288
rect 694 264 699 266
rect 694 262 695 264
rect 697 262 699 264
rect 694 257 699 262
rect 694 255 695 257
rect 697 255 699 257
rect 694 253 699 255
rect 605 250 606 252
rect 608 250 610 252
rect 605 248 610 250
rect 686 252 699 253
rect 686 250 687 252
rect 689 250 699 252
rect 686 249 699 250
rect -1 239 703 243
rect -1 99 3 239
rect 14 231 703 239
rect 11 230 705 231
rect 11 228 31 230
rect 33 228 375 230
rect 377 228 705 230
rect 11 227 705 228
rect 18 221 30 222
rect 18 219 20 221
rect 22 219 30 221
rect 18 216 30 219
rect 18 214 22 216
rect 18 212 20 214
rect 18 189 22 212
rect 130 220 143 221
rect 130 218 140 220
rect 142 218 143 220
rect 130 217 143 218
rect 231 217 244 221
rect 362 221 374 222
rect 333 217 346 221
rect 42 212 64 214
rect 138 215 143 217
rect 138 213 139 215
rect 141 213 143 215
rect 42 210 61 212
rect 63 210 64 212
rect 42 208 54 210
rect 18 187 23 189
rect 18 185 20 187
rect 22 185 23 187
rect 18 180 23 185
rect 34 198 38 206
rect 34 196 46 198
rect 34 194 37 196
rect 39 195 46 196
rect 39 194 40 195
rect 34 193 40 194
rect 42 193 46 195
rect 34 192 46 193
rect 50 196 54 208
rect 52 194 54 196
rect 50 192 54 194
rect 58 205 64 210
rect 58 203 61 205
rect 63 203 64 205
rect 58 201 64 203
rect 18 178 20 180
rect 22 178 23 180
rect 18 176 23 178
rect 58 181 62 201
rect 74 204 112 205
rect 74 202 109 204
rect 111 202 112 204
rect 74 201 112 202
rect 107 198 112 201
rect 82 196 97 197
rect 82 194 86 196
rect 88 194 93 196
rect 95 194 97 196
rect 82 193 97 194
rect 107 196 115 198
rect 107 194 112 196
rect 114 194 115 196
rect 91 187 95 193
rect 107 192 115 194
rect 138 208 143 213
rect 138 206 139 208
rect 141 206 143 208
rect 138 204 143 206
rect 91 185 92 187
rect 94 185 95 187
rect 91 184 95 185
rect 58 180 80 181
rect 58 178 61 180
rect 63 178 80 180
rect 58 177 80 178
rect 139 182 143 204
rect 138 180 143 182
rect 138 178 139 180
rect 141 178 143 180
rect 138 176 143 178
rect 159 212 165 214
rect 239 215 244 217
rect 239 213 240 215
rect 242 213 244 215
rect 159 210 162 212
rect 164 210 165 212
rect 159 205 165 210
rect 159 203 162 205
rect 164 203 165 205
rect 159 201 165 203
rect 159 181 163 201
rect 175 204 213 205
rect 175 202 197 204
rect 199 202 213 204
rect 175 201 213 202
rect 208 198 213 201
rect 183 196 198 197
rect 183 194 187 196
rect 189 194 194 196
rect 196 194 198 196
rect 183 193 198 194
rect 208 196 216 198
rect 208 194 213 196
rect 215 194 216 196
rect 192 184 196 193
rect 208 192 216 194
rect 239 208 244 213
rect 239 206 240 208
rect 242 206 244 208
rect 239 204 244 206
rect 159 180 181 181
rect 159 178 162 180
rect 164 178 181 180
rect 159 177 181 178
rect 240 182 244 204
rect 239 180 244 182
rect 239 178 240 180
rect 242 178 244 180
rect 239 176 244 178
rect 261 212 267 214
rect 341 215 346 217
rect 341 213 342 215
rect 344 213 346 215
rect 261 210 264 212
rect 266 210 267 212
rect 261 205 267 210
rect 261 203 264 205
rect 266 203 267 205
rect 261 201 267 203
rect 261 181 265 201
rect 277 204 315 205
rect 277 202 278 204
rect 280 202 315 204
rect 277 201 315 202
rect 310 198 315 201
rect 285 196 300 197
rect 285 194 289 196
rect 291 194 296 196
rect 298 194 300 196
rect 285 193 300 194
rect 310 196 318 198
rect 310 194 315 196
rect 317 194 318 196
rect 294 187 298 193
rect 310 192 318 194
rect 341 208 346 213
rect 341 206 342 208
rect 344 206 346 208
rect 341 204 346 206
rect 294 185 295 187
rect 297 185 298 187
rect 294 184 298 185
rect 261 180 283 181
rect 261 178 264 180
rect 266 178 283 180
rect 261 177 283 178
rect 342 182 346 204
rect 341 180 346 182
rect 341 178 342 180
rect 344 178 346 180
rect 341 176 346 178
rect 362 219 364 221
rect 366 219 374 221
rect 362 216 374 219
rect 362 214 366 216
rect 362 212 364 214
rect 362 196 366 212
rect 486 217 499 221
rect 587 217 600 221
rect 686 217 699 221
rect 362 194 363 196
rect 365 194 366 196
rect 362 189 366 194
rect 386 212 420 214
rect 494 215 499 217
rect 494 213 495 215
rect 497 213 499 215
rect 386 210 417 212
rect 419 210 420 212
rect 386 208 398 210
rect 362 187 367 189
rect 362 185 364 187
rect 366 185 367 187
rect 362 180 367 185
rect 378 198 382 206
rect 378 196 390 198
rect 378 194 381 196
rect 383 195 390 196
rect 383 194 386 195
rect 378 193 386 194
rect 388 193 390 195
rect 378 192 390 193
rect 394 196 398 208
rect 396 194 398 196
rect 394 192 398 194
rect 414 205 420 210
rect 414 203 417 205
rect 419 203 420 205
rect 414 201 420 203
rect 362 178 364 180
rect 366 178 367 180
rect 362 176 367 178
rect 414 181 418 201
rect 430 204 468 205
rect 430 202 431 204
rect 433 202 468 204
rect 430 201 468 202
rect 463 198 468 201
rect 438 196 453 197
rect 438 194 442 196
rect 444 194 449 196
rect 451 194 453 196
rect 438 193 453 194
rect 463 196 471 198
rect 463 194 468 196
rect 470 194 471 196
rect 447 184 451 193
rect 463 192 471 194
rect 494 208 499 213
rect 494 206 495 208
rect 497 206 499 208
rect 494 204 499 206
rect 414 180 436 181
rect 414 178 417 180
rect 419 178 436 180
rect 414 177 436 178
rect 495 182 499 204
rect 494 180 499 182
rect 491 179 495 180
rect 491 177 492 179
rect 494 178 495 179
rect 497 178 499 180
rect 494 177 499 178
rect 515 212 521 214
rect 595 215 600 217
rect 595 213 596 215
rect 598 213 600 215
rect 515 210 518 212
rect 520 210 521 212
rect 515 205 521 210
rect 515 203 518 205
rect 520 203 521 205
rect 515 201 521 203
rect 515 187 519 201
rect 531 204 569 205
rect 531 202 532 204
rect 534 202 569 204
rect 531 201 569 202
rect 564 198 569 201
rect 539 196 554 197
rect 539 194 543 196
rect 545 194 550 196
rect 552 194 554 196
rect 539 193 554 194
rect 564 196 572 198
rect 564 194 569 196
rect 571 194 572 196
rect 515 185 516 187
rect 518 185 519 187
rect 515 181 519 185
rect 548 187 552 193
rect 564 192 572 194
rect 595 208 600 213
rect 595 206 596 208
rect 598 206 600 208
rect 595 204 600 206
rect 596 195 600 204
rect 596 193 597 195
rect 599 193 600 195
rect 548 185 549 187
rect 551 185 552 187
rect 548 184 552 185
rect 515 180 537 181
rect 515 178 518 180
rect 520 178 537 180
rect 515 177 537 178
rect 596 182 600 193
rect 595 180 600 182
rect 595 178 596 180
rect 598 178 600 180
rect 491 176 499 177
rect 595 176 600 178
rect 614 212 620 214
rect 694 215 699 217
rect 694 213 695 215
rect 697 213 699 215
rect 614 210 617 212
rect 619 210 620 212
rect 614 205 620 210
rect 614 203 617 205
rect 619 203 620 205
rect 614 201 620 203
rect 614 187 618 201
rect 630 204 668 205
rect 630 202 631 204
rect 633 202 668 204
rect 630 201 668 202
rect 663 198 668 201
rect 638 196 653 197
rect 638 194 639 196
rect 641 194 642 196
rect 644 194 649 196
rect 651 194 653 196
rect 638 193 653 194
rect 663 196 671 198
rect 663 194 668 196
rect 670 194 671 196
rect 614 185 615 187
rect 617 185 618 187
rect 614 181 618 185
rect 647 184 651 193
rect 663 192 671 194
rect 694 208 699 213
rect 694 206 695 208
rect 697 206 699 208
rect 694 204 699 206
rect 614 180 636 181
rect 614 178 617 180
rect 619 178 636 180
rect 614 177 636 178
rect 695 182 699 204
rect 694 180 699 182
rect 694 178 695 180
rect 697 178 699 180
rect 694 176 699 178
rect 711 171 715 299
rect 14 170 715 171
rect 14 168 391 170
rect 393 168 715 170
rect 14 167 715 168
rect 14 159 703 167
rect 11 158 703 159
rect 11 156 137 158
rect 139 156 391 158
rect 393 156 703 158
rect 11 155 703 156
rect 19 148 41 149
rect 19 146 22 148
rect 24 146 38 148
rect 40 146 41 148
rect 19 145 41 146
rect 99 148 104 150
rect 99 146 100 148
rect 102 146 104 148
rect 19 125 23 145
rect 52 140 56 142
rect 52 138 53 140
rect 55 138 56 140
rect 19 123 25 125
rect 19 121 22 123
rect 24 121 25 123
rect 19 116 25 121
rect 19 114 22 116
rect 24 114 25 116
rect 19 112 25 114
rect 52 133 56 138
rect 99 144 104 146
rect 43 132 58 133
rect 43 130 47 132
rect 49 130 54 132
rect 56 130 58 132
rect 43 129 58 130
rect 68 132 76 134
rect 68 130 73 132
rect 75 130 76 132
rect 68 128 76 130
rect 68 125 73 128
rect 35 124 73 125
rect 35 122 70 124
rect 72 122 73 124
rect 35 121 73 122
rect 100 122 104 144
rect 99 120 104 122
rect 99 118 100 120
rect 102 118 104 120
rect 99 113 104 118
rect 99 111 100 113
rect 102 111 104 113
rect 99 109 104 111
rect 91 105 104 109
rect 108 148 113 150
rect 108 146 110 148
rect 112 146 113 148
rect 108 141 113 146
rect 160 148 182 149
rect 160 146 163 148
rect 165 146 182 148
rect 160 145 182 146
rect 240 148 245 150
rect 240 146 241 148
rect 243 146 245 148
rect 108 139 110 141
rect 112 139 113 141
rect 108 137 113 139
rect 108 114 112 137
rect 160 134 164 145
rect 193 141 197 142
rect 193 139 194 141
rect 196 139 197 141
rect 124 133 136 134
rect 124 132 132 133
rect 124 130 127 132
rect 129 131 132 132
rect 134 131 136 133
rect 129 130 136 131
rect 124 128 136 130
rect 124 120 128 128
rect 140 132 164 134
rect 142 130 164 132
rect 140 118 144 130
rect 108 112 110 114
rect 108 110 112 112
rect 108 107 120 110
rect 108 105 110 107
rect 112 105 120 107
rect 108 104 120 105
rect 132 112 144 118
rect 160 125 164 130
rect 160 123 166 125
rect 160 121 163 123
rect 165 121 166 123
rect 160 116 166 121
rect 160 114 163 116
rect 165 114 166 116
rect 160 112 166 114
rect 193 133 197 139
rect 240 144 245 146
rect 241 140 245 144
rect 241 138 242 140
rect 244 138 245 140
rect 184 132 199 133
rect 184 130 188 132
rect 190 130 195 132
rect 197 130 199 132
rect 184 129 199 130
rect 209 132 217 134
rect 209 130 214 132
rect 216 130 217 132
rect 209 128 217 130
rect 209 125 214 128
rect 176 121 214 125
rect 241 122 245 138
rect 240 120 245 122
rect 240 118 241 120
rect 243 118 245 120
rect 240 113 245 118
rect 240 111 241 113
rect 243 111 245 113
rect 240 109 245 111
rect 232 105 245 109
rect 261 148 266 150
rect 261 146 263 148
rect 265 146 266 148
rect 261 144 266 146
rect 261 122 265 144
rect 324 148 346 149
rect 324 146 325 148
rect 327 146 341 148
rect 343 146 346 148
rect 324 145 346 146
rect 309 140 313 142
rect 309 138 310 140
rect 312 138 313 140
rect 261 120 266 122
rect 261 118 263 120
rect 265 118 266 120
rect 261 113 266 118
rect 289 132 297 134
rect 309 133 313 138
rect 289 130 290 132
rect 292 130 297 132
rect 289 128 297 130
rect 307 132 322 133
rect 307 130 309 132
rect 311 130 316 132
rect 318 130 322 132
rect 307 129 322 130
rect 292 125 297 128
rect 292 124 330 125
rect 292 122 327 124
rect 329 122 330 124
rect 292 121 330 122
rect 342 125 346 145
rect 340 123 346 125
rect 340 121 341 123
rect 343 121 346 123
rect 340 116 346 121
rect 340 114 341 116
rect 343 114 346 116
rect 261 111 263 113
rect 265 111 266 113
rect 261 109 266 111
rect 340 112 346 114
rect 362 148 367 150
rect 362 146 364 148
rect 366 146 367 148
rect 362 141 367 146
rect 414 148 436 149
rect 414 146 417 148
rect 419 146 436 148
rect 414 145 436 146
rect 494 148 499 150
rect 494 146 495 148
rect 497 146 499 148
rect 362 139 364 141
rect 366 139 367 141
rect 362 137 367 139
rect 362 124 366 137
rect 362 122 363 124
rect 365 122 366 124
rect 362 114 366 122
rect 378 133 390 134
rect 378 132 386 133
rect 378 130 381 132
rect 383 131 386 132
rect 388 131 390 133
rect 383 130 390 131
rect 378 128 390 130
rect 378 120 382 128
rect 394 132 398 134
rect 396 130 398 132
rect 394 118 398 130
rect 362 112 364 114
rect 362 110 366 112
rect 261 108 274 109
rect 261 106 271 108
rect 273 106 274 108
rect 261 105 274 106
rect 362 107 374 110
rect 362 105 364 107
rect 366 105 374 107
rect 362 104 374 105
rect 386 116 398 118
rect 414 125 418 145
rect 414 123 420 125
rect 414 121 417 123
rect 419 121 420 123
rect 414 116 420 121
rect 386 114 417 116
rect 419 114 420 116
rect 386 112 420 114
rect 447 133 451 142
rect 494 144 499 146
rect 438 132 453 133
rect 438 130 442 132
rect 444 130 449 132
rect 451 130 453 132
rect 438 129 453 130
rect 463 132 471 134
rect 463 130 468 132
rect 470 130 471 132
rect 463 128 471 130
rect 463 125 468 128
rect 430 124 468 125
rect 430 122 465 124
rect 467 122 468 124
rect 430 121 468 122
rect 495 122 499 144
rect 494 120 499 122
rect 494 118 495 120
rect 497 118 499 120
rect 494 113 499 118
rect 494 111 495 113
rect 497 111 499 113
rect 515 148 537 149
rect 515 146 518 148
rect 520 146 537 148
rect 515 145 537 146
rect 595 148 600 150
rect 595 146 596 148
rect 598 146 600 148
rect 515 141 519 145
rect 515 139 516 141
rect 518 139 519 141
rect 515 125 519 139
rect 548 141 552 142
rect 548 139 549 141
rect 551 139 552 141
rect 515 123 521 125
rect 515 121 518 123
rect 520 121 521 123
rect 515 116 521 121
rect 515 114 518 116
rect 520 114 521 116
rect 515 112 521 114
rect 548 133 552 139
rect 595 144 600 146
rect 539 132 554 133
rect 539 130 543 132
rect 545 130 550 132
rect 552 130 554 132
rect 539 129 554 130
rect 564 132 572 134
rect 564 130 569 132
rect 571 130 572 132
rect 564 128 572 130
rect 564 125 569 128
rect 596 133 600 144
rect 596 131 597 133
rect 599 131 600 133
rect 531 123 566 125
rect 568 123 569 125
rect 531 121 569 123
rect 596 122 600 131
rect 595 120 600 122
rect 595 118 596 120
rect 598 118 600 120
rect 595 113 600 118
rect 494 109 499 111
rect 595 111 596 113
rect 598 111 600 113
rect 614 148 636 149
rect 614 146 617 148
rect 619 146 636 148
rect 614 145 636 146
rect 694 148 699 150
rect 694 146 695 148
rect 697 146 699 148
rect 614 141 618 145
rect 614 139 615 141
rect 617 139 618 141
rect 614 125 618 139
rect 647 141 651 142
rect 647 139 648 141
rect 650 139 651 141
rect 614 123 620 125
rect 614 121 617 123
rect 619 121 620 123
rect 614 116 620 121
rect 614 114 617 116
rect 619 114 620 116
rect 614 112 620 114
rect 647 133 651 139
rect 694 144 699 146
rect 638 132 653 133
rect 638 130 642 132
rect 644 130 649 132
rect 651 130 653 132
rect 638 129 653 130
rect 663 132 671 134
rect 663 130 668 132
rect 670 130 671 132
rect 663 128 671 130
rect 663 125 668 128
rect 630 124 668 125
rect 630 122 665 124
rect 667 122 668 124
rect 630 121 668 122
rect 695 122 699 144
rect 694 120 699 122
rect 694 118 695 120
rect 697 118 699 120
rect 694 113 699 118
rect 595 109 600 111
rect 694 111 695 113
rect 697 111 699 113
rect 694 109 699 111
rect 486 105 499 109
rect 587 105 600 109
rect 686 105 699 109
rect -1 98 705 99
rect -1 96 121 98
rect 123 96 375 98
rect 377 96 705 98
rect -1 95 705 96
rect -1 94 703 95
rect 11 91 703 94
rect 14 86 702 91
rect 14 84 31 86
rect 33 84 374 86
rect 376 84 702 86
rect 14 83 702 84
rect 18 77 30 78
rect 18 75 20 77
rect 22 75 30 77
rect 18 72 30 75
rect 18 70 22 72
rect 18 68 20 70
rect 18 45 22 68
rect 130 73 143 77
rect 231 73 244 77
rect 361 77 373 78
rect 332 73 345 77
rect 42 68 64 70
rect 138 71 143 73
rect 138 69 139 71
rect 141 69 143 71
rect 42 66 61 68
rect 63 66 64 68
rect 42 64 54 66
rect 18 43 23 45
rect 18 41 20 43
rect 22 41 23 43
rect 18 36 23 41
rect 34 54 38 62
rect 34 52 46 54
rect 34 50 37 52
rect 39 51 46 52
rect 39 50 42 51
rect 34 49 42 50
rect 44 49 46 51
rect 34 48 46 49
rect 50 52 54 64
rect 52 50 54 52
rect 50 48 54 50
rect 58 61 64 66
rect 58 59 61 61
rect 63 59 64 61
rect 58 57 64 59
rect 18 34 20 36
rect 22 34 23 36
rect 18 32 23 34
rect 58 37 62 57
rect 74 60 112 61
rect 74 58 75 60
rect 77 58 112 60
rect 74 57 112 58
rect 107 54 112 57
rect 82 52 97 53
rect 82 50 86 52
rect 88 50 93 52
rect 95 50 97 52
rect 82 49 97 50
rect 107 52 115 54
rect 107 50 112 52
rect 114 50 115 52
rect 91 40 95 49
rect 107 48 115 50
rect 138 64 143 69
rect 138 62 139 64
rect 141 62 143 64
rect 138 60 143 62
rect 58 36 80 37
rect 58 34 61 36
rect 63 34 80 36
rect 58 33 80 34
rect 139 38 143 60
rect 138 36 143 38
rect 138 34 139 36
rect 141 34 143 36
rect 138 32 143 34
rect 159 68 165 70
rect 239 71 244 73
rect 239 69 240 71
rect 242 69 244 71
rect 159 66 162 68
rect 164 66 165 68
rect 159 61 165 66
rect 159 59 162 61
rect 164 59 165 61
rect 159 57 165 59
rect 159 43 163 57
rect 175 60 213 61
rect 175 58 176 60
rect 178 58 213 60
rect 175 57 213 58
rect 208 54 213 57
rect 183 52 198 53
rect 183 50 187 52
rect 189 50 194 52
rect 196 50 198 52
rect 183 49 198 50
rect 208 52 216 54
rect 208 50 213 52
rect 215 50 216 52
rect 159 41 160 43
rect 162 41 163 43
rect 159 37 163 41
rect 192 43 196 49
rect 208 48 216 50
rect 239 64 244 69
rect 239 62 240 64
rect 242 62 244 64
rect 239 60 244 62
rect 240 51 244 60
rect 240 49 241 51
rect 243 49 244 51
rect 192 41 193 43
rect 195 41 196 43
rect 192 40 196 41
rect 159 36 181 37
rect 159 34 162 36
rect 164 34 181 36
rect 159 33 181 34
rect 240 38 244 49
rect 239 36 244 38
rect 239 34 240 36
rect 242 34 244 36
rect 239 32 244 34
rect 260 68 266 70
rect 340 71 345 73
rect 340 69 341 71
rect 343 69 345 71
rect 260 66 263 68
rect 265 66 266 68
rect 260 61 266 66
rect 260 59 263 61
rect 265 59 266 61
rect 260 57 266 59
rect 260 43 264 57
rect 276 60 314 61
rect 276 58 277 60
rect 279 58 314 60
rect 276 57 314 58
rect 309 54 314 57
rect 284 52 299 53
rect 284 50 288 52
rect 290 50 295 52
rect 297 50 299 52
rect 284 49 299 50
rect 309 52 317 54
rect 309 50 314 52
rect 316 50 317 52
rect 293 48 297 49
rect 309 48 317 50
rect 260 41 261 43
rect 263 41 264 43
rect 293 46 294 48
rect 296 46 297 48
rect 260 37 264 41
rect 293 40 297 46
rect 340 64 345 69
rect 340 62 341 64
rect 343 62 345 64
rect 340 60 345 62
rect 260 36 282 37
rect 260 34 263 36
rect 265 34 282 36
rect 260 33 282 34
rect 341 38 345 60
rect 340 36 345 38
rect 340 34 341 36
rect 343 34 345 36
rect 340 32 345 34
rect 361 75 363 77
rect 365 75 373 77
rect 361 72 373 75
rect 361 70 365 72
rect 361 68 363 70
rect 361 48 365 68
rect 485 73 498 77
rect 586 73 599 77
rect 685 73 698 77
rect 361 46 362 48
rect 364 46 365 48
rect 361 45 365 46
rect 385 68 419 70
rect 493 71 498 73
rect 493 69 494 71
rect 496 69 498 71
rect 385 66 416 68
rect 418 66 419 68
rect 385 64 397 66
rect 361 43 366 45
rect 361 41 363 43
rect 365 41 366 43
rect 361 36 366 41
rect 377 54 381 62
rect 377 52 389 54
rect 377 50 380 52
rect 382 51 389 52
rect 382 50 385 51
rect 377 49 385 50
rect 387 49 389 51
rect 377 48 389 49
rect 393 52 397 64
rect 395 50 397 52
rect 393 48 397 50
rect 413 61 419 66
rect 413 59 416 61
rect 418 59 419 61
rect 413 57 419 59
rect 361 34 363 36
rect 365 34 366 36
rect 361 32 366 34
rect 413 37 417 57
rect 429 60 467 61
rect 429 58 430 60
rect 432 58 467 60
rect 429 57 467 58
rect 462 54 467 57
rect 437 52 452 53
rect 437 50 441 52
rect 443 50 448 52
rect 450 50 452 52
rect 437 49 452 50
rect 462 52 470 54
rect 462 50 467 52
rect 469 50 470 52
rect 446 40 450 49
rect 462 48 470 50
rect 493 64 498 69
rect 493 62 494 64
rect 496 62 498 64
rect 493 60 498 62
rect 413 36 435 37
rect 413 34 416 36
rect 418 34 435 36
rect 413 33 435 34
rect 494 38 498 60
rect 493 36 498 38
rect 493 34 494 36
rect 496 34 498 36
rect 493 32 498 34
rect 514 68 520 70
rect 594 71 599 73
rect 594 69 595 71
rect 597 69 599 71
rect 514 66 517 68
rect 519 66 520 68
rect 514 61 520 66
rect 514 59 517 61
rect 519 59 520 61
rect 514 57 520 59
rect 514 43 518 57
rect 530 60 568 61
rect 530 58 531 60
rect 533 58 568 60
rect 530 57 568 58
rect 563 54 568 57
rect 538 52 553 53
rect 538 50 542 52
rect 544 50 549 52
rect 551 50 553 52
rect 538 49 553 50
rect 563 52 571 54
rect 563 50 568 52
rect 570 50 571 52
rect 514 41 515 43
rect 517 41 518 43
rect 514 37 518 41
rect 547 43 551 49
rect 563 48 571 50
rect 594 64 599 69
rect 594 62 595 64
rect 597 62 599 64
rect 594 60 599 62
rect 595 51 599 60
rect 595 49 596 51
rect 598 49 599 51
rect 547 41 548 43
rect 550 41 551 43
rect 547 40 551 41
rect 514 36 536 37
rect 514 34 517 36
rect 519 34 536 36
rect 514 33 536 34
rect 595 38 599 49
rect 594 36 599 38
rect 594 34 595 36
rect 597 34 599 36
rect 594 32 599 34
rect 613 68 619 70
rect 693 71 698 73
rect 693 69 694 71
rect 696 69 698 71
rect 613 66 616 68
rect 618 66 619 68
rect 613 61 619 66
rect 613 59 616 61
rect 618 59 619 61
rect 613 57 619 59
rect 613 43 617 57
rect 629 60 667 61
rect 629 58 630 60
rect 632 58 667 60
rect 629 57 667 58
rect 662 54 667 57
rect 637 52 652 53
rect 637 50 638 52
rect 640 50 641 52
rect 643 50 648 52
rect 650 50 652 52
rect 637 49 652 50
rect 662 52 670 54
rect 662 50 667 52
rect 669 50 670 52
rect 613 41 614 43
rect 616 41 617 43
rect 613 37 617 41
rect 646 40 650 49
rect 662 48 670 50
rect 693 64 698 69
rect 693 62 694 64
rect 696 62 698 64
rect 693 60 698 62
rect 613 36 635 37
rect 613 34 616 36
rect 618 34 635 36
rect 613 33 635 34
rect 694 38 698 60
rect 693 36 698 38
rect 693 34 694 36
rect 696 34 698 36
rect 693 32 698 34
rect 711 27 715 167
rect 11 26 715 27
rect 11 24 47 26
rect 49 24 390 26
rect 392 24 715 26
rect 11 23 715 24
rect 14 19 702 23
<< alu2 >>
rect 347 372 547 373
rect 347 370 348 372
rect 350 370 544 372
rect 546 370 547 372
rect 347 369 547 370
rect 49 364 118 365
rect 49 362 50 364
rect 52 362 115 364
rect 117 362 118 364
rect 49 361 118 362
rect 260 364 329 365
rect 260 362 261 364
rect 263 362 326 364
rect 328 362 329 364
rect 260 361 329 362
rect 430 364 499 365
rect 430 362 431 364
rect 433 362 496 364
rect 498 362 499 364
rect 430 361 499 362
rect 565 364 634 365
rect 565 362 566 364
rect 568 362 631 364
rect 633 362 634 364
rect 565 361 634 362
rect 58 356 490 357
rect 58 354 59 356
rect 61 354 487 356
rect 489 354 490 356
rect 58 353 490 354
rect 27 348 62 349
rect 27 346 28 348
rect 30 346 59 348
rect 61 346 62 348
rect 27 345 62 346
rect 114 348 118 349
rect 114 346 115 348
rect 117 346 118 348
rect 114 345 118 346
rect 260 348 264 349
rect 260 346 261 348
rect 263 346 264 348
rect 260 345 264 346
rect 316 348 351 349
rect 316 346 317 348
rect 319 346 348 348
rect 350 346 351 348
rect 316 345 351 346
rect 430 348 434 349
rect 430 346 431 348
rect 433 346 434 348
rect 430 345 434 346
rect 486 348 521 349
rect 486 346 487 348
rect 489 346 518 348
rect 520 346 521 348
rect 486 345 521 346
rect 543 348 578 349
rect 543 346 544 348
rect 546 346 575 348
rect 577 346 578 348
rect 543 345 578 346
rect 630 348 634 349
rect 630 346 631 348
rect 633 346 634 348
rect 630 345 634 346
rect 25 340 353 341
rect 25 338 26 340
rect 28 338 350 340
rect 352 338 353 340
rect 25 337 353 338
rect 479 339 585 340
rect 479 337 480 339
rect 482 337 582 339
rect 584 337 585 339
rect 479 336 585 337
rect 25 331 29 332
rect 25 329 26 331
rect 28 329 29 331
rect 25 328 29 329
rect 65 331 69 332
rect 65 329 66 331
rect 68 329 69 331
rect 65 328 69 329
rect 131 331 135 332
rect 131 329 132 331
rect 134 329 135 331
rect 131 328 135 329
rect 243 331 247 332
rect 243 329 244 331
rect 246 329 247 331
rect 243 328 247 329
rect 309 331 313 332
rect 309 329 310 331
rect 312 329 313 331
rect 309 328 313 329
rect 349 331 353 332
rect 349 329 350 331
rect 352 329 353 331
rect 349 328 353 329
rect 413 331 417 332
rect 413 329 414 331
rect 416 329 417 331
rect 413 328 417 329
rect 479 331 483 332
rect 479 329 480 331
rect 482 329 483 331
rect 479 328 483 329
rect 519 331 523 332
rect 519 329 520 331
rect 522 329 523 331
rect 519 328 523 329
rect 541 331 545 332
rect 541 329 542 331
rect 544 329 545 331
rect 541 328 545 329
rect 581 331 585 332
rect 581 329 582 331
rect 584 329 585 331
rect 581 328 585 329
rect 647 331 651 332
rect 647 329 648 331
rect 650 329 651 331
rect 647 328 651 329
rect 116 324 120 325
rect 89 323 97 324
rect 89 321 90 323
rect 92 321 94 323
rect 96 321 97 323
rect 116 322 117 324
rect 119 322 120 324
rect 116 321 120 322
rect 178 324 187 325
rect 178 322 179 324
rect 181 322 184 324
rect 186 322 187 324
rect 178 321 187 322
rect 196 324 200 325
rect 196 322 197 324
rect 199 322 200 324
rect 196 321 200 322
rect 258 324 262 325
rect 366 324 370 325
rect 258 322 259 324
rect 261 322 262 324
rect 258 321 262 322
rect 281 323 289 324
rect 281 321 282 323
rect 284 321 286 323
rect 288 321 289 323
rect 366 322 367 324
rect 369 322 370 324
rect 366 321 370 322
rect 428 324 432 325
rect 632 324 636 325
rect 428 322 429 324
rect 431 322 432 324
rect 428 321 432 322
rect 451 323 459 324
rect 451 321 452 323
rect 454 321 456 323
rect 458 321 459 323
rect 89 320 97 321
rect 281 320 289 321
rect 451 320 459 321
rect 605 323 613 324
rect 605 321 606 323
rect 608 321 610 323
rect 612 321 613 323
rect 632 322 633 324
rect 635 322 636 324
rect 632 321 636 322
rect 605 320 613 321
rect 89 293 135 294
rect 89 291 90 293
rect 92 291 132 293
rect 134 291 135 293
rect 89 290 135 291
rect 243 293 289 294
rect 243 291 244 293
rect 246 291 286 293
rect 288 291 289 293
rect 243 290 289 291
rect 413 293 459 294
rect 413 291 414 293
rect 416 291 456 293
rect 458 291 459 293
rect 413 290 459 291
rect 605 293 651 294
rect 605 291 606 293
rect 608 291 648 293
rect 650 291 651 293
rect 605 290 651 291
rect 25 285 29 286
rect 25 283 26 285
rect 28 283 29 285
rect 25 282 29 283
rect 65 285 313 286
rect 65 283 66 285
rect 68 283 310 285
rect 312 283 313 285
rect 65 282 313 283
rect 349 285 353 286
rect 479 285 483 286
rect 349 283 350 285
rect 352 283 353 285
rect 349 282 353 283
rect 405 284 450 285
rect 405 282 406 284
rect 408 282 447 284
rect 449 282 450 284
rect 479 283 480 285
rect 482 283 483 285
rect 479 282 483 283
rect 519 285 545 286
rect 519 283 520 285
rect 522 283 542 285
rect 544 283 545 285
rect 519 282 545 283
rect 581 285 585 286
rect 581 283 582 285
rect 584 283 585 285
rect 581 282 585 283
rect 405 281 450 282
rect 46 276 54 277
rect 46 274 47 276
rect 49 274 51 276
rect 53 274 54 276
rect 46 273 54 274
rect 116 276 126 277
rect 116 274 117 276
rect 119 274 123 276
rect 125 274 126 276
rect 116 273 126 274
rect 195 276 248 277
rect 195 274 196 276
rect 198 274 245 276
rect 247 274 248 276
rect 195 273 248 274
rect 252 276 262 277
rect 252 274 253 276
rect 255 274 259 276
rect 261 274 262 276
rect 252 273 262 274
rect 422 276 432 277
rect 422 274 423 276
rect 425 274 429 276
rect 431 274 432 276
rect 422 273 432 274
rect 494 276 509 277
rect 494 274 495 276
rect 497 274 506 276
rect 508 274 509 276
rect 494 273 509 274
rect 632 276 642 277
rect 632 274 633 276
rect 635 274 639 276
rect 641 274 642 276
rect 632 273 642 274
rect 27 268 62 269
rect 27 266 28 268
rect 30 266 55 268
rect 57 266 59 268
rect 61 266 62 268
rect 27 265 62 266
rect 93 268 118 269
rect 93 266 94 268
rect 96 266 115 268
rect 117 266 118 268
rect 93 265 118 266
rect 155 268 209 269
rect 155 266 156 268
rect 158 266 206 268
rect 208 266 209 268
rect 155 265 209 266
rect 260 268 285 269
rect 260 266 261 268
rect 263 266 282 268
rect 284 266 285 268
rect 260 265 285 266
rect 316 268 351 269
rect 316 266 317 268
rect 319 266 348 268
rect 350 266 351 268
rect 316 265 351 266
rect 430 268 455 269
rect 430 266 431 268
rect 433 266 452 268
rect 454 266 455 268
rect 430 265 455 266
rect 486 268 521 269
rect 486 266 487 268
rect 489 266 518 268
rect 520 266 521 268
rect 486 265 521 266
rect 543 268 578 269
rect 543 266 544 268
rect 546 266 575 268
rect 577 266 578 268
rect 543 265 578 266
rect 609 268 634 269
rect 609 266 610 268
rect 612 266 631 268
rect 633 266 634 268
rect 609 265 634 266
rect 356 264 370 265
rect 356 262 357 264
rect 359 262 367 264
rect 369 262 370 264
rect 356 261 370 262
rect 100 260 104 261
rect 100 258 101 260
rect 103 258 104 260
rect 205 260 278 261
rect 205 258 206 260
rect 208 258 275 260
rect 277 258 278 260
rect 100 257 104 258
rect 174 257 182 258
rect 174 255 175 257
rect 177 255 179 257
rect 181 255 182 257
rect 174 254 182 255
rect 196 257 200 258
rect 205 257 278 258
rect 600 260 620 261
rect 600 258 601 260
rect 603 258 617 260
rect 619 258 620 260
rect 600 257 620 258
rect 196 255 197 257
rect 199 255 200 257
rect 196 254 200 255
rect 325 255 329 256
rect 325 253 326 255
rect 328 253 329 255
rect 325 252 329 253
rect 347 255 547 256
rect 347 253 348 255
rect 350 253 544 255
rect 546 253 547 255
rect 347 252 547 253
rect 686 252 690 253
rect 686 250 687 252
rect 689 250 690 252
rect 686 249 690 250
rect 54 247 490 248
rect 54 245 55 247
rect 57 245 487 247
rect 489 245 490 247
rect 54 244 490 245
rect 139 220 281 221
rect 139 218 140 220
rect 142 218 278 220
rect 280 218 281 220
rect 139 217 281 218
rect 325 220 634 221
rect 325 218 326 220
rect 328 218 631 220
rect 633 218 634 220
rect 325 217 634 218
rect 244 212 434 213
rect 244 210 245 212
rect 247 210 431 212
rect 433 210 434 212
rect 244 209 434 210
rect 505 212 642 213
rect 505 210 506 212
rect 508 210 639 212
rect 641 210 642 212
rect 505 209 642 210
rect 108 204 151 205
rect 108 202 109 204
rect 111 202 148 204
rect 150 202 151 204
rect 108 201 151 202
rect 196 204 200 205
rect 196 202 197 204
rect 199 202 200 204
rect 196 201 200 202
rect 277 204 281 205
rect 277 202 278 204
rect 280 202 281 204
rect 277 201 281 202
rect 305 204 409 205
rect 305 202 306 204
rect 308 202 406 204
rect 408 202 409 204
rect 305 201 409 202
rect 430 204 434 205
rect 430 202 431 204
rect 433 202 434 204
rect 430 201 434 202
rect 531 204 535 205
rect 531 202 532 204
rect 534 202 535 204
rect 531 201 535 202
rect 630 204 634 205
rect 630 202 631 204
rect 633 202 634 204
rect 630 201 634 202
rect 193 196 366 197
rect 448 196 452 197
rect 638 196 642 197
rect 39 195 43 196
rect 39 193 40 195
rect 42 193 43 195
rect 39 192 43 193
rect 100 195 112 196
rect 100 193 101 195
rect 103 193 109 195
rect 111 193 112 195
rect 193 194 194 196
rect 196 194 363 196
rect 365 194 366 196
rect 193 193 366 194
rect 385 195 389 196
rect 385 193 386 195
rect 388 193 389 195
rect 100 192 112 193
rect 147 188 255 189
rect 385 188 389 193
rect 448 194 449 196
rect 451 195 600 196
rect 451 194 597 195
rect 448 193 597 194
rect 599 193 600 195
rect 638 194 639 196
rect 641 194 642 196
rect 638 193 642 194
rect 448 192 600 193
rect 91 187 103 188
rect 91 185 92 187
rect 94 185 100 187
rect 102 185 103 187
rect 147 186 148 188
rect 150 186 252 188
rect 254 186 255 188
rect 147 185 255 186
rect 294 187 298 188
rect 294 185 295 187
rect 297 185 298 187
rect 91 184 103 185
rect 294 184 298 185
rect 385 187 519 188
rect 385 185 516 187
rect 518 185 519 187
rect 385 184 519 185
rect 548 187 618 188
rect 548 185 549 187
rect 551 185 615 187
rect 617 185 618 187
rect 548 184 618 185
rect 19 180 23 181
rect 19 178 20 180
rect 22 178 23 180
rect 19 177 23 178
rect 131 180 165 181
rect 131 178 132 180
rect 134 178 162 180
rect 164 178 165 180
rect 131 177 165 178
rect 192 180 243 181
rect 341 180 345 181
rect 647 180 698 181
rect 192 178 194 180
rect 196 178 240 180
rect 242 178 243 180
rect 192 177 243 178
rect 251 179 309 180
rect 251 177 252 179
rect 254 177 306 179
rect 308 177 309 179
rect 341 178 342 180
rect 344 178 345 180
rect 341 177 345 178
rect 491 179 495 180
rect 491 177 492 179
rect 494 177 495 179
rect 647 178 648 180
rect 650 178 695 180
rect 697 178 698 180
rect 647 177 698 178
rect 251 176 309 177
rect 491 176 495 177
rect 366 171 535 172
rect 366 169 367 171
rect 369 169 532 171
rect 534 169 535 171
rect 366 168 535 169
rect 37 148 41 149
rect 37 146 38 148
rect 40 146 41 148
rect 37 145 41 146
rect 99 148 103 149
rect 99 146 100 148
rect 102 146 103 148
rect 99 145 103 146
rect 294 148 328 149
rect 294 146 295 148
rect 297 146 325 148
rect 327 146 328 148
rect 294 145 328 146
rect 109 141 113 142
rect 52 140 110 141
rect 52 138 53 140
rect 55 139 110 140
rect 112 139 113 141
rect 55 138 113 139
rect 193 141 197 142
rect 385 141 519 142
rect 193 139 194 141
rect 196 139 197 141
rect 193 138 197 139
rect 241 140 313 141
rect 241 138 242 140
rect 244 138 310 140
rect 312 138 313 140
rect 52 137 113 138
rect 241 137 313 138
rect 385 139 516 141
rect 518 139 519 141
rect 385 138 519 139
rect 548 141 618 142
rect 548 139 549 141
rect 551 139 615 141
rect 617 139 618 141
rect 548 138 618 139
rect 647 141 651 142
rect 647 139 648 141
rect 650 139 651 141
rect 647 138 651 139
rect 131 133 135 134
rect 385 133 389 138
rect 131 131 132 133
rect 134 131 135 133
rect 131 130 135 131
rect 213 132 360 133
rect 213 130 214 132
rect 216 130 357 132
rect 359 130 360 132
rect 385 131 386 133
rect 388 131 389 133
rect 385 130 389 131
rect 448 133 600 134
rect 448 132 597 133
rect 448 130 449 132
rect 451 131 597 132
rect 599 131 600 133
rect 451 130 600 131
rect 213 129 360 130
rect 448 129 452 130
rect 565 125 604 126
rect 69 124 159 125
rect 69 122 70 124
rect 72 122 156 124
rect 158 122 159 124
rect 69 121 159 122
rect 326 124 366 125
rect 326 122 327 124
rect 329 122 363 124
rect 365 122 366 124
rect 326 121 366 122
rect 464 124 495 125
rect 464 122 465 124
rect 467 122 492 124
rect 494 122 495 124
rect 565 123 566 125
rect 568 123 601 125
rect 603 123 604 125
rect 565 122 604 123
rect 664 124 690 125
rect 664 122 665 124
rect 667 122 687 124
rect 689 122 690 124
rect 464 121 495 122
rect 664 121 690 122
rect 270 108 274 109
rect 270 106 271 108
rect 273 106 274 108
rect 270 105 274 106
rect 270 100 641 101
rect 270 98 271 100
rect 273 98 638 100
rect 640 98 641 100
rect 270 97 641 98
rect 341 82 433 83
rect 341 80 342 82
rect 344 80 430 82
rect 432 80 433 82
rect 341 79 433 80
rect 174 68 280 69
rect 174 66 175 68
rect 177 66 277 68
rect 279 66 280 68
rect 174 65 280 66
rect 19 60 78 61
rect 19 58 20 60
rect 22 58 75 60
rect 77 58 78 60
rect 19 57 78 58
rect 108 60 179 61
rect 108 58 109 60
rect 111 58 176 60
rect 178 58 179 60
rect 108 57 179 58
rect 276 60 280 61
rect 276 58 277 60
rect 279 58 280 60
rect 276 57 280 58
rect 429 60 433 61
rect 429 58 430 60
rect 432 58 433 60
rect 429 57 433 58
rect 530 60 534 61
rect 530 58 531 60
rect 533 58 534 60
rect 530 57 534 58
rect 629 60 633 61
rect 629 58 630 60
rect 632 58 633 60
rect 629 57 633 58
rect 92 52 96 53
rect 447 52 451 53
rect 637 52 641 53
rect 41 51 45 52
rect 41 49 42 51
rect 44 49 45 51
rect 41 44 45 49
rect 92 50 93 52
rect 95 51 244 52
rect 95 50 241 51
rect 92 49 241 50
rect 243 49 244 51
rect 384 51 388 52
rect 384 49 385 51
rect 387 49 388 51
rect 92 48 244 49
rect 293 48 365 49
rect 293 46 294 48
rect 296 46 362 48
rect 364 46 365 48
rect 293 45 365 46
rect 384 44 388 49
rect 447 50 448 52
rect 450 51 599 52
rect 450 50 596 51
rect 447 49 596 50
rect 598 49 599 51
rect 637 50 638 52
rect 640 50 641 52
rect 637 49 641 50
rect 447 48 599 49
rect 41 43 163 44
rect 41 41 160 43
rect 162 41 163 43
rect 41 40 163 41
rect 192 43 264 44
rect 192 41 193 43
rect 195 41 261 43
rect 263 41 264 43
rect 192 40 264 41
rect 384 43 518 44
rect 384 41 515 43
rect 517 41 518 43
rect 384 40 518 41
rect 547 43 617 44
rect 547 41 548 43
rect 550 41 614 43
rect 616 41 617 43
rect 547 40 617 41
rect 183 35 534 36
rect 183 33 184 35
rect 186 33 531 35
rect 533 33 534 35
rect 183 32 534 33
rect 47 27 633 28
rect 47 25 48 27
rect 50 25 630 27
rect 632 25 633 27
rect 47 24 633 25
<< alu3 >>
rect 347 372 351 373
rect 347 370 348 372
rect 350 370 351 372
rect 114 364 118 365
rect 114 362 115 364
rect 117 362 118 364
rect 58 356 62 357
rect 58 354 59 356
rect 61 354 62 356
rect 58 348 62 354
rect 58 346 59 348
rect 61 346 62 348
rect 58 345 62 346
rect 114 348 118 362
rect 114 346 115 348
rect 117 346 118 348
rect 114 345 118 346
rect 260 364 264 365
rect 260 362 261 364
rect 263 362 264 364
rect 260 348 264 362
rect 260 346 261 348
rect 263 346 264 348
rect 260 345 264 346
rect 347 348 351 370
rect 543 372 547 373
rect 543 370 544 372
rect 546 370 547 372
rect 347 346 348 348
rect 350 346 351 348
rect 347 345 351 346
rect 430 364 434 365
rect 430 362 431 364
rect 433 362 434 364
rect 430 348 434 362
rect 430 346 431 348
rect 433 346 434 348
rect 430 345 434 346
rect 486 356 490 357
rect 486 354 487 356
rect 489 354 490 356
rect 486 348 490 354
rect 486 346 487 348
rect 489 346 490 348
rect 486 345 490 346
rect 543 348 547 370
rect 543 346 544 348
rect 546 346 547 348
rect 543 345 547 346
rect 630 364 634 365
rect 630 362 631 364
rect 633 362 634 364
rect 630 348 634 362
rect 630 346 631 348
rect 633 346 634 348
rect 630 345 634 346
rect 25 340 29 341
rect 25 338 26 340
rect 28 338 29 340
rect 25 331 29 338
rect 349 340 353 341
rect 349 338 350 340
rect 352 338 353 340
rect 25 329 26 331
rect 28 329 29 331
rect 25 285 29 329
rect 25 283 26 285
rect 28 283 29 285
rect 25 282 29 283
rect 65 331 69 332
rect 65 329 66 331
rect 68 329 69 331
rect 65 285 69 329
rect 131 331 135 332
rect 131 329 132 331
rect 134 329 135 331
rect 116 324 120 325
rect 65 283 66 285
rect 68 283 69 285
rect 65 282 69 283
rect 93 323 97 324
rect 93 321 94 323
rect 96 321 97 323
rect 46 276 50 277
rect 46 274 47 276
rect 49 274 50 276
rect 46 204 50 274
rect 54 268 58 269
rect 54 266 55 268
rect 57 266 58 268
rect 54 247 58 266
rect 93 268 97 321
rect 116 322 117 324
rect 119 322 120 324
rect 116 276 120 322
rect 131 293 135 329
rect 243 331 247 332
rect 243 329 244 331
rect 246 329 247 331
rect 131 291 132 293
rect 134 291 135 293
rect 131 290 135 291
rect 183 324 187 325
rect 183 322 184 324
rect 186 322 187 324
rect 116 274 117 276
rect 119 274 120 276
rect 116 273 120 274
rect 93 266 94 268
rect 96 266 97 268
rect 93 265 97 266
rect 155 268 159 269
rect 155 266 156 268
rect 158 266 159 268
rect 54 245 55 247
rect 57 245 58 247
rect 54 244 58 245
rect 100 260 104 261
rect 100 258 101 260
rect 103 258 104 260
rect 46 200 51 204
rect 37 195 43 196
rect 37 193 40 195
rect 42 193 43 195
rect 37 192 43 193
rect 19 180 23 181
rect 19 178 20 180
rect 22 178 23 180
rect 19 60 23 178
rect 37 148 41 192
rect 37 146 38 148
rect 40 146 41 148
rect 37 145 41 146
rect 19 58 20 60
rect 22 58 23 60
rect 19 57 23 58
rect 47 27 51 200
rect 100 195 104 258
rect 147 204 151 205
rect 147 202 148 204
rect 150 202 151 204
rect 100 193 101 195
rect 103 193 104 195
rect 100 192 104 193
rect 108 195 112 196
rect 108 193 109 195
rect 111 193 112 195
rect 99 187 103 188
rect 99 185 100 187
rect 102 185 103 187
rect 99 148 103 185
rect 99 146 100 148
rect 102 146 103 148
rect 99 145 103 146
rect 108 60 112 193
rect 147 188 151 202
rect 147 186 148 188
rect 150 186 151 188
rect 147 185 151 186
rect 131 180 135 181
rect 131 178 132 180
rect 134 178 135 180
rect 131 133 135 178
rect 131 131 132 133
rect 134 131 135 133
rect 131 130 135 131
rect 155 124 159 266
rect 155 122 156 124
rect 158 122 159 124
rect 155 121 159 122
rect 174 257 178 258
rect 174 255 175 257
rect 177 255 178 257
rect 174 68 178 255
rect 174 66 175 68
rect 177 66 178 68
rect 174 65 178 66
rect 108 58 109 60
rect 111 58 112 60
rect 108 57 112 58
rect 183 35 187 322
rect 195 324 200 325
rect 195 322 197 324
rect 199 322 200 324
rect 195 321 200 322
rect 195 276 199 321
rect 243 293 247 329
rect 309 331 313 332
rect 309 329 310 331
rect 312 329 313 331
rect 243 291 244 293
rect 246 291 247 293
rect 243 290 247 291
rect 258 324 262 325
rect 258 322 259 324
rect 261 322 262 324
rect 195 274 196 276
rect 198 274 199 276
rect 195 273 199 274
rect 244 276 248 277
rect 244 274 245 276
rect 247 274 248 276
rect 205 268 209 269
rect 205 266 206 268
rect 208 266 209 268
rect 205 260 209 266
rect 205 258 206 260
rect 208 258 209 260
rect 196 257 200 258
rect 205 257 209 258
rect 196 255 197 257
rect 199 255 200 257
rect 196 204 200 255
rect 244 212 248 274
rect 258 276 262 322
rect 258 274 259 276
rect 261 274 262 276
rect 258 273 262 274
rect 281 323 285 324
rect 281 321 282 323
rect 284 321 285 323
rect 281 268 285 321
rect 309 285 313 329
rect 309 283 310 285
rect 312 283 313 285
rect 309 282 313 283
rect 349 331 353 338
rect 479 339 483 340
rect 479 337 480 339
rect 482 337 483 339
rect 349 329 350 331
rect 352 329 353 331
rect 349 285 353 329
rect 413 331 417 332
rect 413 329 414 331
rect 416 329 417 331
rect 349 283 350 285
rect 352 283 353 285
rect 349 282 353 283
rect 366 324 370 325
rect 366 322 367 324
rect 369 322 370 324
rect 281 266 282 268
rect 284 266 285 268
rect 281 265 285 266
rect 347 268 351 269
rect 347 266 348 268
rect 350 266 351 268
rect 325 255 329 256
rect 325 253 326 255
rect 328 253 329 255
rect 244 210 245 212
rect 247 210 248 212
rect 244 209 248 210
rect 277 220 281 221
rect 277 218 278 220
rect 280 218 281 220
rect 196 202 197 204
rect 199 202 200 204
rect 196 201 200 202
rect 277 204 281 218
rect 325 220 329 253
rect 347 255 351 266
rect 347 253 348 255
rect 350 253 351 255
rect 347 252 351 253
rect 356 264 360 265
rect 356 262 357 264
rect 359 262 360 264
rect 325 218 326 220
rect 328 218 329 220
rect 325 217 329 218
rect 277 202 278 204
rect 280 202 281 204
rect 277 201 281 202
rect 305 204 309 205
rect 305 202 306 204
rect 308 202 309 204
rect 251 188 255 189
rect 251 186 252 188
rect 254 186 255 188
rect 193 180 197 181
rect 193 178 194 180
rect 196 178 197 180
rect 193 141 197 178
rect 251 179 255 186
rect 251 177 252 179
rect 254 177 255 179
rect 251 176 255 177
rect 294 187 298 188
rect 294 185 295 187
rect 297 185 298 187
rect 294 148 298 185
rect 305 179 309 202
rect 305 177 306 179
rect 308 177 309 179
rect 305 176 309 177
rect 341 180 345 181
rect 341 178 342 180
rect 344 178 345 180
rect 294 146 295 148
rect 297 146 298 148
rect 294 145 298 146
rect 193 139 194 141
rect 196 139 197 141
rect 193 138 197 139
rect 270 108 274 109
rect 270 106 271 108
rect 273 106 274 108
rect 270 100 274 106
rect 270 98 271 100
rect 273 98 274 100
rect 270 97 274 98
rect 341 82 345 178
rect 356 132 360 262
rect 366 171 370 322
rect 413 293 417 329
rect 479 331 483 337
rect 581 339 585 340
rect 581 337 582 339
rect 584 337 585 339
rect 479 329 480 331
rect 482 329 483 331
rect 413 291 414 293
rect 416 291 417 293
rect 413 290 417 291
rect 428 324 432 325
rect 428 322 429 324
rect 431 322 432 324
rect 405 284 409 285
rect 405 282 406 284
rect 408 282 409 284
rect 405 204 409 282
rect 428 276 432 322
rect 428 274 429 276
rect 431 274 432 276
rect 428 273 432 274
rect 451 323 455 324
rect 451 321 452 323
rect 454 321 455 323
rect 451 268 455 321
rect 479 285 483 329
rect 479 283 480 285
rect 482 283 483 285
rect 479 282 483 283
rect 519 331 523 332
rect 519 329 520 331
rect 522 329 523 331
rect 519 285 523 329
rect 519 283 520 285
rect 522 283 523 285
rect 519 282 523 283
rect 541 331 545 332
rect 541 329 542 331
rect 544 329 545 331
rect 541 285 545 329
rect 541 283 542 285
rect 544 283 545 285
rect 541 282 545 283
rect 581 331 585 337
rect 581 329 582 331
rect 584 329 585 331
rect 581 285 585 329
rect 647 331 651 332
rect 647 329 648 331
rect 650 329 651 331
rect 632 324 636 325
rect 581 283 582 285
rect 584 283 585 285
rect 581 282 585 283
rect 609 323 613 324
rect 609 321 610 323
rect 612 321 613 323
rect 505 276 509 277
rect 505 274 506 276
rect 508 274 509 276
rect 451 266 452 268
rect 454 266 455 268
rect 451 265 455 266
rect 486 268 490 269
rect 486 266 487 268
rect 489 266 490 268
rect 486 247 490 266
rect 486 245 487 247
rect 489 245 490 247
rect 486 244 490 245
rect 405 202 406 204
rect 408 202 409 204
rect 405 201 409 202
rect 430 212 434 213
rect 430 210 431 212
rect 433 210 434 212
rect 430 204 434 210
rect 505 212 509 274
rect 543 268 547 269
rect 543 266 544 268
rect 546 266 547 268
rect 543 255 547 266
rect 609 268 613 321
rect 632 322 633 324
rect 635 322 636 324
rect 632 276 636 322
rect 647 293 651 329
rect 647 291 648 293
rect 650 291 651 293
rect 647 290 651 291
rect 632 274 633 276
rect 635 274 636 276
rect 632 273 636 274
rect 609 266 610 268
rect 612 266 613 268
rect 609 265 613 266
rect 543 253 544 255
rect 546 253 547 255
rect 543 252 547 253
rect 600 260 604 261
rect 600 258 601 260
rect 603 258 604 260
rect 505 210 506 212
rect 508 210 509 212
rect 505 209 509 210
rect 430 202 431 204
rect 433 202 434 204
rect 430 201 434 202
rect 531 204 535 205
rect 531 202 532 204
rect 534 202 535 204
rect 366 169 367 171
rect 369 169 370 171
rect 366 168 370 169
rect 491 179 495 180
rect 491 177 492 179
rect 494 177 495 179
rect 356 130 357 132
rect 359 130 360 132
rect 356 129 360 130
rect 491 124 495 177
rect 531 171 535 202
rect 531 169 532 171
rect 534 169 535 171
rect 531 168 535 169
rect 491 122 492 124
rect 494 122 495 124
rect 600 125 604 258
rect 686 252 690 253
rect 686 250 687 252
rect 689 250 690 252
rect 630 220 634 221
rect 630 218 631 220
rect 633 218 634 220
rect 630 204 634 218
rect 630 202 631 204
rect 633 202 634 204
rect 630 201 634 202
rect 638 212 642 213
rect 638 210 639 212
rect 641 210 642 212
rect 638 196 642 210
rect 638 194 639 196
rect 641 194 642 196
rect 638 193 642 194
rect 647 180 651 181
rect 647 178 648 180
rect 650 178 651 180
rect 647 141 651 178
rect 647 139 648 141
rect 650 139 651 141
rect 647 138 651 139
rect 600 123 601 125
rect 603 123 604 125
rect 600 122 604 123
rect 686 124 690 250
rect 686 122 687 124
rect 689 122 690 124
rect 491 121 495 122
rect 686 121 690 122
rect 637 100 641 101
rect 637 98 638 100
rect 640 98 641 100
rect 341 80 342 82
rect 344 80 345 82
rect 341 79 345 80
rect 429 82 433 83
rect 429 80 430 82
rect 432 80 433 82
rect 276 68 280 69
rect 276 66 277 68
rect 279 66 280 68
rect 276 60 280 66
rect 276 58 277 60
rect 279 58 280 60
rect 276 57 280 58
rect 429 60 433 80
rect 429 58 430 60
rect 432 58 433 60
rect 429 57 433 58
rect 530 60 534 61
rect 530 58 531 60
rect 533 58 534 60
rect 183 33 184 35
rect 186 33 187 35
rect 183 32 187 33
rect 530 35 534 58
rect 530 33 531 35
rect 533 33 534 35
rect 530 32 534 33
rect 629 60 633 61
rect 629 58 630 60
rect 632 58 633 60
rect 47 25 48 27
rect 50 25 51 27
rect 47 24 51 25
rect 629 27 633 58
rect 637 52 641 98
rect 637 50 638 52
rect 640 50 641 52
rect 637 49 641 50
rect 629 25 630 27
rect 632 25 633 27
rect 629 24 633 25
<< ptie >>
rect 43 166 53 172
rect 387 170 397 172
rect 387 168 391 170
rect 393 168 397 170
rect 387 166 397 168
rect 133 158 143 160
rect 133 156 137 158
rect 139 156 143 158
rect 133 154 143 156
rect 387 158 397 160
rect 387 156 391 158
rect 393 156 397 158
rect 387 154 397 156
rect 43 26 53 28
rect 43 24 47 26
rect 49 24 53 26
rect 43 22 53 24
rect 386 26 396 28
rect 386 24 390 26
rect 392 24 396 26
rect 386 22 396 24
<< nmos >>
rect 25 320 27 333
rect 32 320 34 333
rect 45 319 47 333
rect 65 320 67 333
rect 72 320 74 333
rect 85 319 87 333
rect 106 313 108 327
rect 117 313 119 333
rect 124 313 126 333
rect 144 319 146 333
rect 154 319 156 333
rect 164 316 166 326
rect 174 313 176 326
rect 202 313 204 326
rect 212 316 214 326
rect 222 319 224 333
rect 232 319 234 333
rect 252 313 254 333
rect 259 313 261 333
rect 270 313 272 327
rect 291 319 293 333
rect 304 320 306 333
rect 311 320 313 333
rect 331 319 333 333
rect 344 320 346 333
rect 351 320 353 333
rect 372 313 374 326
rect 382 316 384 326
rect 392 319 394 333
rect 402 319 404 333
rect 422 313 424 333
rect 429 313 431 333
rect 440 313 442 327
rect 461 319 463 333
rect 474 320 476 333
rect 481 320 483 333
rect 501 319 503 333
rect 514 320 516 333
rect 521 320 523 333
rect 541 320 543 333
rect 548 320 550 333
rect 561 319 563 333
rect 581 320 583 333
rect 588 320 590 333
rect 601 319 603 333
rect 622 313 624 327
rect 633 313 635 333
rect 640 313 642 333
rect 660 319 662 333
rect 670 319 672 333
rect 680 316 682 326
rect 690 313 692 326
rect 25 281 27 294
rect 32 281 34 294
rect 45 281 47 295
rect 65 281 67 294
rect 72 281 74 294
rect 85 281 87 295
rect 106 287 108 301
rect 117 281 119 301
rect 124 281 126 301
rect 144 281 146 295
rect 154 281 156 295
rect 164 288 166 298
rect 174 288 176 301
rect 202 288 204 301
rect 212 288 214 298
rect 222 281 224 295
rect 232 281 234 295
rect 252 281 254 301
rect 259 281 261 301
rect 270 287 272 301
rect 291 281 293 295
rect 304 281 306 294
rect 311 281 313 294
rect 331 281 333 295
rect 344 281 346 294
rect 351 281 353 294
rect 372 288 374 301
rect 382 288 384 298
rect 392 281 394 295
rect 402 281 404 295
rect 422 281 424 301
rect 429 281 431 301
rect 440 287 442 301
rect 461 281 463 295
rect 474 281 476 294
rect 481 281 483 294
rect 501 281 503 295
rect 514 281 516 294
rect 521 281 523 294
rect 541 281 543 294
rect 548 281 550 294
rect 561 281 563 295
rect 581 281 583 294
rect 588 281 590 294
rect 601 281 603 295
rect 622 287 624 301
rect 633 281 635 301
rect 640 281 642 301
rect 660 281 662 295
rect 670 281 672 295
rect 680 288 682 298
rect 690 288 692 301
rect 25 175 27 189
rect 35 176 37 184
rect 45 178 47 186
rect 66 169 68 183
rect 77 169 79 189
rect 84 169 86 189
rect 104 175 106 189
rect 114 175 116 189
rect 124 172 126 182
rect 134 169 136 182
rect 167 169 169 183
rect 178 169 180 189
rect 185 169 187 189
rect 205 175 207 189
rect 215 175 217 189
rect 225 172 227 182
rect 235 169 237 182
rect 269 169 271 183
rect 280 169 282 189
rect 287 169 289 189
rect 307 175 309 189
rect 317 175 319 189
rect 327 172 329 182
rect 337 169 339 182
rect 369 175 371 189
rect 379 176 381 184
rect 389 178 391 186
rect 422 169 424 183
rect 433 169 435 189
rect 440 169 442 189
rect 460 175 462 189
rect 470 175 472 189
rect 480 172 482 182
rect 490 169 492 182
rect 523 169 525 183
rect 534 169 536 189
rect 541 169 543 189
rect 561 175 563 189
rect 571 175 573 189
rect 581 172 583 182
rect 591 169 593 182
rect 622 169 624 183
rect 633 169 635 189
rect 640 169 642 189
rect 660 175 662 189
rect 670 175 672 189
rect 680 172 682 182
rect 690 169 692 182
rect 27 143 29 157
rect 38 137 40 157
rect 45 137 47 157
rect 65 137 67 151
rect 75 137 77 151
rect 85 144 87 154
rect 95 144 97 157
rect 115 137 117 151
rect 125 142 127 150
rect 135 140 137 148
rect 168 143 170 157
rect 179 137 181 157
rect 186 137 188 157
rect 206 137 208 151
rect 216 137 218 151
rect 226 144 228 154
rect 236 144 238 157
rect 268 144 270 157
rect 278 144 280 154
rect 288 137 290 151
rect 298 137 300 151
rect 318 137 320 157
rect 325 137 327 157
rect 336 143 338 157
rect 369 137 371 151
rect 379 142 381 150
rect 389 140 391 148
rect 422 143 424 157
rect 433 137 435 157
rect 440 137 442 157
rect 460 137 462 151
rect 470 137 472 151
rect 480 144 482 154
rect 490 144 492 157
rect 523 143 525 157
rect 534 137 536 157
rect 541 137 543 157
rect 561 137 563 151
rect 571 137 573 151
rect 581 144 583 154
rect 591 144 593 157
rect 622 143 624 157
rect 633 137 635 157
rect 640 137 642 157
rect 660 137 662 151
rect 670 137 672 151
rect 680 144 682 154
rect 690 144 692 157
rect 25 31 27 45
rect 35 32 37 40
rect 45 34 47 42
rect 66 25 68 39
rect 77 25 79 45
rect 84 25 86 45
rect 104 31 106 45
rect 114 31 116 45
rect 124 28 126 38
rect 134 25 136 38
rect 167 25 169 39
rect 178 25 180 45
rect 185 25 187 45
rect 205 31 207 45
rect 215 31 217 45
rect 225 28 227 38
rect 235 25 237 38
rect 268 25 270 39
rect 279 25 281 45
rect 286 25 288 45
rect 306 31 308 45
rect 316 31 318 45
rect 326 28 328 38
rect 336 25 338 38
rect 368 31 370 45
rect 378 32 380 40
rect 388 34 390 42
rect 421 25 423 39
rect 432 25 434 45
rect 439 25 441 45
rect 459 31 461 45
rect 469 31 471 45
rect 479 28 481 38
rect 489 25 491 38
rect 522 25 524 39
rect 533 25 535 45
rect 540 25 542 45
rect 560 31 562 45
rect 570 31 572 45
rect 580 28 582 38
rect 590 25 592 38
rect 621 25 623 39
rect 632 25 634 45
rect 639 25 641 45
rect 659 31 661 45
rect 669 31 671 45
rect 679 28 681 38
rect 689 25 691 38
<< pmos >>
rect 25 354 27 373
rect 35 354 37 373
rect 45 345 47 373
rect 65 354 67 373
rect 75 354 77 373
rect 85 345 87 373
rect 106 345 108 373
rect 116 345 118 373
rect 126 345 128 373
rect 144 345 146 370
rect 151 345 153 370
rect 161 348 163 361
rect 174 348 176 373
rect 202 348 204 373
rect 215 348 217 361
rect 225 345 227 370
rect 232 345 234 370
rect 250 345 252 373
rect 260 345 262 373
rect 270 345 272 373
rect 291 345 293 373
rect 301 354 303 373
rect 311 354 313 373
rect 331 345 333 373
rect 341 354 343 373
rect 351 354 353 373
rect 372 348 374 373
rect 385 348 387 361
rect 395 345 397 370
rect 402 345 404 370
rect 420 345 422 373
rect 430 345 432 373
rect 440 345 442 373
rect 461 345 463 373
rect 471 354 473 373
rect 481 354 483 373
rect 501 345 503 373
rect 511 354 513 373
rect 521 354 523 373
rect 541 354 543 373
rect 551 354 553 373
rect 561 345 563 373
rect 581 354 583 373
rect 591 354 593 373
rect 601 345 603 373
rect 622 345 624 373
rect 632 345 634 373
rect 642 345 644 373
rect 660 345 662 370
rect 667 345 669 370
rect 677 348 679 361
rect 690 348 692 373
rect 25 241 27 260
rect 35 241 37 260
rect 45 241 47 269
rect 65 241 67 260
rect 75 241 77 260
rect 85 241 87 269
rect 106 241 108 269
rect 116 241 118 269
rect 126 241 128 269
rect 144 244 146 269
rect 151 244 153 269
rect 161 253 163 266
rect 174 241 176 266
rect 202 241 204 266
rect 215 253 217 266
rect 225 244 227 269
rect 232 244 234 269
rect 250 241 252 269
rect 260 241 262 269
rect 270 241 272 269
rect 291 241 293 269
rect 301 241 303 260
rect 311 241 313 260
rect 331 241 333 269
rect 341 241 343 260
rect 351 241 353 260
rect 372 241 374 266
rect 385 253 387 266
rect 395 244 397 269
rect 402 244 404 269
rect 420 241 422 269
rect 430 241 432 269
rect 440 241 442 269
rect 461 241 463 269
rect 471 241 473 260
rect 481 241 483 260
rect 501 241 503 269
rect 511 241 513 260
rect 521 241 523 260
rect 541 241 543 260
rect 551 241 553 260
rect 561 241 563 269
rect 581 241 583 260
rect 591 241 593 260
rect 601 241 603 269
rect 622 241 624 269
rect 632 241 634 269
rect 642 241 644 269
rect 660 244 662 269
rect 667 244 669 269
rect 677 253 679 266
rect 690 241 692 266
rect 25 201 27 229
rect 38 201 40 229
rect 45 201 47 229
rect 66 201 68 229
rect 76 201 78 229
rect 86 201 88 229
rect 104 201 106 226
rect 111 201 113 226
rect 121 204 123 217
rect 134 204 136 229
rect 167 201 169 229
rect 177 201 179 229
rect 187 201 189 229
rect 205 201 207 226
rect 212 201 214 226
rect 222 204 224 217
rect 235 204 237 229
rect 269 201 271 229
rect 279 201 281 229
rect 289 201 291 229
rect 307 201 309 226
rect 314 201 316 226
rect 324 204 326 217
rect 337 204 339 229
rect 369 201 371 229
rect 382 201 384 229
rect 389 201 391 229
rect 422 201 424 229
rect 432 201 434 229
rect 442 201 444 229
rect 460 201 462 226
rect 467 201 469 226
rect 477 204 479 217
rect 490 204 492 229
rect 523 201 525 229
rect 533 201 535 229
rect 543 201 545 229
rect 561 201 563 226
rect 568 201 570 226
rect 578 204 580 217
rect 591 204 593 229
rect 622 201 624 229
rect 632 201 634 229
rect 642 201 644 229
rect 660 201 662 226
rect 667 201 669 226
rect 677 204 679 217
rect 690 204 692 229
rect 27 97 29 125
rect 37 97 39 125
rect 47 97 49 125
rect 65 100 67 125
rect 72 100 74 125
rect 82 109 84 122
rect 95 97 97 122
rect 115 97 117 125
rect 128 97 130 125
rect 135 97 137 125
rect 168 97 170 125
rect 178 97 180 125
rect 188 97 190 125
rect 206 100 208 125
rect 213 100 215 125
rect 223 109 225 122
rect 236 97 238 122
rect 268 97 270 122
rect 281 109 283 122
rect 291 100 293 125
rect 298 100 300 125
rect 316 97 318 125
rect 326 97 328 125
rect 336 97 338 125
rect 369 97 371 125
rect 382 97 384 125
rect 389 97 391 125
rect 422 97 424 125
rect 432 97 434 125
rect 442 97 444 125
rect 460 100 462 125
rect 467 100 469 125
rect 477 109 479 122
rect 490 97 492 122
rect 523 97 525 125
rect 533 97 535 125
rect 543 97 545 125
rect 561 100 563 125
rect 568 100 570 125
rect 578 109 580 122
rect 591 97 593 122
rect 622 97 624 125
rect 632 97 634 125
rect 642 97 644 125
rect 660 100 662 125
rect 667 100 669 125
rect 677 109 679 122
rect 690 97 692 122
rect 25 57 27 85
rect 38 57 40 85
rect 45 57 47 85
rect 66 57 68 85
rect 76 57 78 85
rect 86 57 88 85
rect 104 57 106 82
rect 111 57 113 82
rect 121 60 123 73
rect 134 60 136 85
rect 167 57 169 85
rect 177 57 179 85
rect 187 57 189 85
rect 205 57 207 82
rect 212 57 214 82
rect 222 60 224 73
rect 235 60 237 85
rect 268 57 270 85
rect 278 57 280 85
rect 288 57 290 85
rect 306 57 308 82
rect 313 57 315 82
rect 323 60 325 73
rect 336 60 338 85
rect 368 57 370 85
rect 381 57 383 85
rect 388 57 390 85
rect 421 57 423 85
rect 431 57 433 85
rect 441 57 443 85
rect 459 57 461 82
rect 466 57 468 82
rect 476 60 478 73
rect 489 60 491 85
rect 522 57 524 85
rect 532 57 534 85
rect 542 57 544 85
rect 560 57 562 82
rect 567 57 569 82
rect 577 60 579 73
rect 590 60 592 85
rect 621 57 623 85
rect 631 57 633 85
rect 641 57 643 85
rect 659 57 661 82
rect 666 57 668 82
rect 676 60 678 73
rect 689 60 691 85
<< polyct0 >>
rect 43 338 45 340
rect 83 338 85 340
rect 106 338 108 340
rect 116 338 118 340
rect 166 341 168 343
rect 172 331 174 333
rect 210 341 212 343
rect 204 331 206 333
rect 260 338 262 340
rect 270 338 272 340
rect 293 338 295 340
rect 333 338 335 340
rect 380 341 382 343
rect 374 331 376 333
rect 430 338 432 340
rect 440 338 442 340
rect 463 338 465 340
rect 503 338 505 340
rect 559 338 561 340
rect 599 338 601 340
rect 622 338 624 340
rect 632 338 634 340
rect 682 341 684 343
rect 688 331 690 333
rect 43 274 45 276
rect 83 274 85 276
rect 106 274 108 276
rect 116 274 118 276
rect 172 281 174 283
rect 166 271 168 273
rect 204 281 206 283
rect 210 271 212 273
rect 374 281 376 283
rect 260 274 262 276
rect 270 274 272 276
rect 293 274 295 276
rect 333 274 335 276
rect 380 271 382 273
rect 430 274 432 276
rect 440 274 442 276
rect 463 274 465 276
rect 503 274 505 276
rect 559 274 561 276
rect 599 274 601 276
rect 622 274 624 276
rect 632 274 634 276
rect 688 281 690 283
rect 682 271 684 273
rect 27 194 29 196
rect 66 194 68 196
rect 76 194 78 196
rect 126 197 128 199
rect 167 194 169 196
rect 177 194 179 196
rect 132 187 134 189
rect 227 197 229 199
rect 269 194 271 196
rect 279 194 281 196
rect 233 187 235 189
rect 329 197 331 199
rect 371 194 373 196
rect 422 194 424 196
rect 432 194 434 196
rect 335 187 337 189
rect 482 197 484 199
rect 523 194 525 196
rect 533 194 535 196
rect 488 187 490 189
rect 583 197 585 199
rect 622 194 624 196
rect 632 194 634 196
rect 589 187 591 189
rect 682 197 684 199
rect 688 187 690 189
rect 27 130 29 132
rect 37 130 39 132
rect 93 137 95 139
rect 87 127 89 129
rect 117 130 119 132
rect 168 130 170 132
rect 178 130 180 132
rect 234 137 236 139
rect 228 127 230 129
rect 270 137 272 139
rect 276 127 278 129
rect 326 130 328 132
rect 336 130 338 132
rect 371 130 373 132
rect 422 130 424 132
rect 432 130 434 132
rect 488 137 490 139
rect 482 127 484 129
rect 523 130 525 132
rect 533 130 535 132
rect 589 137 591 139
rect 583 127 585 129
rect 622 130 624 132
rect 632 130 634 132
rect 688 137 690 139
rect 682 127 684 129
rect 27 50 29 52
rect 66 50 68 52
rect 76 50 78 52
rect 126 53 128 55
rect 167 50 169 52
rect 177 50 179 52
rect 132 43 134 45
rect 227 53 229 55
rect 268 50 270 52
rect 278 50 280 52
rect 233 43 235 45
rect 328 53 330 55
rect 370 50 372 52
rect 421 50 423 52
rect 431 50 433 52
rect 334 43 336 45
rect 481 53 483 55
rect 522 50 524 52
rect 532 50 534 52
rect 487 43 489 45
rect 582 53 584 55
rect 621 50 623 52
rect 631 50 633 52
rect 588 43 590 45
rect 681 53 683 55
rect 687 43 689 45
<< polyct1 >>
rect 23 346 25 348
rect 63 346 65 348
rect 33 338 35 340
rect 73 338 75 340
rect 126 338 128 340
rect 133 338 135 340
rect 152 338 154 340
rect 313 346 315 348
rect 224 338 226 340
rect 243 338 245 340
rect 250 338 252 340
rect 303 338 305 340
rect 353 346 355 348
rect 343 338 345 340
rect 483 346 485 348
rect 394 338 396 340
rect 413 338 415 340
rect 420 338 422 340
rect 473 338 475 340
rect 523 346 525 348
rect 539 346 541 348
rect 513 338 515 340
rect 579 346 581 348
rect 549 338 551 340
rect 589 338 591 340
rect 642 338 644 340
rect 649 338 651 340
rect 668 338 670 340
rect 33 274 35 276
rect 23 266 25 268
rect 73 274 75 276
rect 126 274 128 276
rect 133 274 135 276
rect 152 274 154 276
rect 63 266 65 268
rect 224 274 226 276
rect 243 274 245 276
rect 250 274 252 276
rect 303 274 305 276
rect 343 274 345 276
rect 313 266 315 268
rect 353 266 355 268
rect 394 274 396 276
rect 413 274 415 276
rect 420 274 422 276
rect 473 274 475 276
rect 513 274 515 276
rect 483 266 485 268
rect 549 274 551 276
rect 523 266 525 268
rect 539 266 541 268
rect 589 274 591 276
rect 642 274 644 276
rect 649 274 651 276
rect 668 274 670 276
rect 579 266 581 268
rect 37 194 39 196
rect 50 194 52 196
rect 86 194 88 196
rect 93 194 95 196
rect 112 194 114 196
rect 187 194 189 196
rect 194 194 196 196
rect 213 194 215 196
rect 289 194 291 196
rect 296 194 298 196
rect 315 194 317 196
rect 381 194 383 196
rect 394 194 396 196
rect 442 194 444 196
rect 449 194 451 196
rect 468 194 470 196
rect 543 194 545 196
rect 550 194 552 196
rect 569 194 571 196
rect 642 194 644 196
rect 649 194 651 196
rect 668 194 670 196
rect 47 130 49 132
rect 54 130 56 132
rect 73 130 75 132
rect 127 130 129 132
rect 140 130 142 132
rect 188 130 190 132
rect 195 130 197 132
rect 214 130 216 132
rect 290 130 292 132
rect 309 130 311 132
rect 316 130 318 132
rect 381 130 383 132
rect 394 130 396 132
rect 442 130 444 132
rect 449 130 451 132
rect 468 130 470 132
rect 543 130 545 132
rect 550 130 552 132
rect 569 130 571 132
rect 642 130 644 132
rect 649 130 651 132
rect 668 130 670 132
rect 37 50 39 52
rect 50 50 52 52
rect 86 50 88 52
rect 93 50 95 52
rect 112 50 114 52
rect 187 50 189 52
rect 194 50 196 52
rect 213 50 215 52
rect 288 50 290 52
rect 295 50 297 52
rect 314 50 316 52
rect 380 50 382 52
rect 393 50 395 52
rect 441 50 443 52
rect 448 50 450 52
rect 467 50 469 52
rect 542 50 544 52
rect 549 50 551 52
rect 568 50 570 52
rect 641 50 643 52
rect 648 50 650 52
rect 667 50 669 52
<< ndifct0 >>
rect 20 322 22 324
rect 60 322 62 324
rect 112 315 114 317
rect 139 329 141 331
rect 129 322 131 324
rect 139 322 141 324
rect 149 329 151 331
rect 159 321 161 323
rect 169 318 171 320
rect 207 318 209 320
rect 217 321 219 323
rect 227 329 229 331
rect 237 329 239 331
rect 237 322 239 324
rect 247 322 249 324
rect 264 315 266 317
rect 316 322 318 324
rect 356 322 358 324
rect 377 318 379 320
rect 387 321 389 323
rect 397 329 399 331
rect 407 329 409 331
rect 407 322 409 324
rect 417 322 419 324
rect 434 315 436 317
rect 486 322 488 324
rect 526 322 528 324
rect 536 322 538 324
rect 576 322 578 324
rect 628 315 630 317
rect 655 329 657 331
rect 645 322 647 324
rect 655 322 657 324
rect 665 329 667 331
rect 675 321 677 323
rect 685 318 687 320
rect 20 290 22 292
rect 60 290 62 292
rect 112 297 114 299
rect 129 290 131 292
rect 139 290 141 292
rect 139 283 141 285
rect 149 283 151 285
rect 159 291 161 293
rect 169 294 171 296
rect 207 294 209 296
rect 217 291 219 293
rect 227 283 229 285
rect 237 290 239 292
rect 247 290 249 292
rect 237 283 239 285
rect 264 297 266 299
rect 316 290 318 292
rect 356 290 358 292
rect 377 294 379 296
rect 387 291 389 293
rect 397 283 399 285
rect 407 290 409 292
rect 417 290 419 292
rect 407 283 409 285
rect 434 297 436 299
rect 486 290 488 292
rect 526 290 528 292
rect 536 290 538 292
rect 576 290 578 292
rect 628 297 630 299
rect 645 290 647 292
rect 655 290 657 292
rect 655 283 657 285
rect 665 283 667 285
rect 675 291 677 293
rect 685 294 687 296
rect 30 178 32 180
rect 40 180 42 182
rect 50 180 52 182
rect 72 171 74 173
rect 99 185 101 187
rect 89 178 91 180
rect 99 178 101 180
rect 109 185 111 187
rect 119 177 121 179
rect 129 174 131 176
rect 173 171 175 173
rect 200 185 202 187
rect 190 178 192 180
rect 200 178 202 180
rect 210 185 212 187
rect 220 177 222 179
rect 230 174 232 176
rect 275 171 277 173
rect 302 185 304 187
rect 292 178 294 180
rect 302 178 304 180
rect 312 185 314 187
rect 322 177 324 179
rect 332 174 334 176
rect 374 178 376 180
rect 384 180 386 182
rect 394 180 396 182
rect 428 171 430 173
rect 455 185 457 187
rect 445 178 447 180
rect 455 178 457 180
rect 465 185 467 187
rect 475 177 477 179
rect 485 174 487 176
rect 529 171 531 173
rect 556 185 558 187
rect 546 178 548 180
rect 556 178 558 180
rect 566 185 568 187
rect 576 177 578 179
rect 586 174 588 176
rect 628 171 630 173
rect 655 185 657 187
rect 645 178 647 180
rect 655 178 657 180
rect 665 185 667 187
rect 675 177 677 179
rect 685 174 687 176
rect 33 153 35 155
rect 50 146 52 148
rect 60 146 62 148
rect 60 139 62 141
rect 70 139 72 141
rect 80 147 82 149
rect 90 150 92 152
rect 120 146 122 148
rect 130 144 132 146
rect 140 144 142 146
rect 174 153 176 155
rect 191 146 193 148
rect 201 146 203 148
rect 201 139 203 141
rect 211 139 213 141
rect 221 147 223 149
rect 231 150 233 152
rect 273 150 275 152
rect 283 147 285 149
rect 293 139 295 141
rect 303 146 305 148
rect 313 146 315 148
rect 303 139 305 141
rect 330 153 332 155
rect 374 146 376 148
rect 384 144 386 146
rect 394 144 396 146
rect 428 153 430 155
rect 445 146 447 148
rect 455 146 457 148
rect 455 139 457 141
rect 465 139 467 141
rect 475 147 477 149
rect 485 150 487 152
rect 529 153 531 155
rect 546 146 548 148
rect 556 146 558 148
rect 556 139 558 141
rect 566 139 568 141
rect 576 147 578 149
rect 586 150 588 152
rect 628 153 630 155
rect 645 146 647 148
rect 655 146 657 148
rect 655 139 657 141
rect 665 139 667 141
rect 675 147 677 149
rect 685 150 687 152
rect 30 34 32 36
rect 40 36 42 38
rect 50 36 52 38
rect 72 27 74 29
rect 99 41 101 43
rect 89 34 91 36
rect 99 34 101 36
rect 109 41 111 43
rect 119 33 121 35
rect 129 30 131 32
rect 173 27 175 29
rect 200 41 202 43
rect 190 34 192 36
rect 200 34 202 36
rect 210 41 212 43
rect 220 33 222 35
rect 230 30 232 32
rect 274 27 276 29
rect 301 41 303 43
rect 291 34 293 36
rect 301 34 303 36
rect 311 41 313 43
rect 321 33 323 35
rect 331 30 333 32
rect 373 34 375 36
rect 383 36 385 38
rect 393 36 395 38
rect 427 27 429 29
rect 454 41 456 43
rect 444 34 446 36
rect 454 34 456 36
rect 464 41 466 43
rect 474 33 476 35
rect 484 30 486 32
rect 528 27 530 29
rect 555 41 557 43
rect 545 34 547 36
rect 555 34 557 36
rect 565 41 567 43
rect 575 33 577 35
rect 585 30 587 32
rect 627 27 629 29
rect 654 41 656 43
rect 644 34 646 36
rect 654 34 656 36
rect 664 41 666 43
rect 674 33 676 35
rect 684 30 686 32
<< ndifct1 >>
rect 50 329 52 331
rect 50 321 52 323
rect 90 329 92 331
rect 90 321 92 323
rect 101 322 103 324
rect 39 312 41 314
rect 79 312 81 314
rect 179 322 181 324
rect 197 322 199 324
rect 286 329 288 331
rect 275 322 277 324
rect 286 321 288 323
rect 326 329 328 331
rect 326 321 328 323
rect 367 322 369 324
rect 297 312 299 314
rect 337 312 339 314
rect 456 329 458 331
rect 445 322 447 324
rect 456 321 458 323
rect 496 329 498 331
rect 496 321 498 323
rect 566 329 568 331
rect 566 321 568 323
rect 467 312 469 314
rect 507 312 509 314
rect 606 329 608 331
rect 606 321 608 323
rect 617 322 619 324
rect 555 312 557 314
rect 595 312 597 314
rect 695 322 697 324
rect 39 300 41 302
rect 79 300 81 302
rect 50 291 52 293
rect 50 283 52 285
rect 90 291 92 293
rect 101 290 103 292
rect 90 283 92 285
rect 179 290 181 292
rect 197 290 199 292
rect 297 300 299 302
rect 337 300 339 302
rect 275 290 277 292
rect 286 291 288 293
rect 286 283 288 285
rect 326 291 328 293
rect 326 283 328 285
rect 367 290 369 292
rect 467 300 469 302
rect 507 300 509 302
rect 445 290 447 292
rect 456 291 458 293
rect 456 283 458 285
rect 555 300 557 302
rect 595 300 597 302
rect 496 291 498 293
rect 496 283 498 285
rect 566 291 568 293
rect 566 283 568 285
rect 606 291 608 293
rect 617 290 619 292
rect 606 283 608 285
rect 695 290 697 292
rect 20 185 22 187
rect 20 178 22 180
rect 61 178 63 180
rect 139 178 141 180
rect 162 178 164 180
rect 240 178 242 180
rect 264 178 266 180
rect 364 185 366 187
rect 342 178 344 180
rect 364 178 366 180
rect 417 178 419 180
rect 495 178 497 180
rect 518 178 520 180
rect 596 178 598 180
rect 617 178 619 180
rect 695 178 697 180
rect 22 146 24 148
rect 100 146 102 148
rect 110 146 112 148
rect 110 139 112 141
rect 163 146 165 148
rect 241 146 243 148
rect 263 146 265 148
rect 341 146 343 148
rect 364 146 366 148
rect 364 139 366 141
rect 417 146 419 148
rect 495 146 497 148
rect 518 146 520 148
rect 596 146 598 148
rect 617 146 619 148
rect 695 146 697 148
rect 20 41 22 43
rect 20 34 22 36
rect 61 34 63 36
rect 139 34 141 36
rect 162 34 164 36
rect 240 34 242 36
rect 263 34 265 36
rect 363 41 365 43
rect 341 34 343 36
rect 363 34 365 36
rect 416 34 418 36
rect 494 34 496 36
rect 517 34 519 36
rect 595 34 597 36
rect 616 34 618 36
rect 694 34 696 36
<< ptiect1 >>
rect 391 168 393 170
rect 137 156 139 158
rect 391 156 393 158
rect 47 24 49 26
rect 390 24 392 26
<< pdifct0 >>
rect 20 369 22 371
rect 20 362 22 364
rect 30 363 32 365
rect 30 356 32 358
rect 40 369 42 371
rect 40 362 42 364
rect 60 369 62 371
rect 60 362 62 364
rect 70 363 72 365
rect 70 356 72 358
rect 80 369 82 371
rect 80 362 82 364
rect 111 369 113 371
rect 111 362 113 364
rect 121 361 123 363
rect 121 354 123 356
rect 133 369 135 371
rect 133 362 135 364
rect 168 369 170 371
rect 156 350 158 352
rect 208 369 210 371
rect 220 350 222 352
rect 243 369 245 371
rect 243 362 245 364
rect 255 361 257 363
rect 255 354 257 356
rect 265 369 267 371
rect 265 362 267 364
rect 296 369 298 371
rect 296 362 298 364
rect 306 363 308 365
rect 306 356 308 358
rect 316 369 318 371
rect 316 362 318 364
rect 336 369 338 371
rect 336 362 338 364
rect 346 363 348 365
rect 346 356 348 358
rect 356 369 358 371
rect 356 362 358 364
rect 378 369 380 371
rect 390 350 392 352
rect 413 369 415 371
rect 413 362 415 364
rect 425 361 427 363
rect 425 354 427 356
rect 435 369 437 371
rect 435 362 437 364
rect 466 369 468 371
rect 466 362 468 364
rect 476 363 478 365
rect 476 356 478 358
rect 486 369 488 371
rect 486 362 488 364
rect 506 369 508 371
rect 506 362 508 364
rect 516 363 518 365
rect 516 356 518 358
rect 526 369 528 371
rect 526 362 528 364
rect 536 369 538 371
rect 536 362 538 364
rect 546 363 548 365
rect 546 356 548 358
rect 556 369 558 371
rect 556 362 558 364
rect 576 369 578 371
rect 576 362 578 364
rect 586 363 588 365
rect 586 356 588 358
rect 596 369 598 371
rect 596 362 598 364
rect 627 369 629 371
rect 627 362 629 364
rect 637 361 639 363
rect 637 354 639 356
rect 649 369 651 371
rect 649 362 651 364
rect 684 369 686 371
rect 672 350 674 352
rect 20 250 22 252
rect 20 243 22 245
rect 30 256 32 258
rect 30 249 32 251
rect 40 250 42 252
rect 40 243 42 245
rect 60 250 62 252
rect 60 243 62 245
rect 70 256 72 258
rect 70 249 72 251
rect 80 250 82 252
rect 80 243 82 245
rect 111 250 113 252
rect 111 243 113 245
rect 121 258 123 260
rect 121 251 123 253
rect 133 250 135 252
rect 133 243 135 245
rect 156 262 158 264
rect 168 243 170 245
rect 220 262 222 264
rect 208 243 210 245
rect 243 250 245 252
rect 243 243 245 245
rect 255 258 257 260
rect 255 251 257 253
rect 265 250 267 252
rect 265 243 267 245
rect 296 250 298 252
rect 296 243 298 245
rect 306 256 308 258
rect 306 249 308 251
rect 316 250 318 252
rect 316 243 318 245
rect 336 250 338 252
rect 336 243 338 245
rect 346 256 348 258
rect 346 249 348 251
rect 356 250 358 252
rect 356 243 358 245
rect 390 262 392 264
rect 378 243 380 245
rect 413 250 415 252
rect 413 243 415 245
rect 425 258 427 260
rect 425 251 427 253
rect 435 250 437 252
rect 435 243 437 245
rect 466 250 468 252
rect 466 243 468 245
rect 476 256 478 258
rect 476 249 478 251
rect 486 250 488 252
rect 486 243 488 245
rect 506 250 508 252
rect 506 243 508 245
rect 516 256 518 258
rect 516 249 518 251
rect 526 250 528 252
rect 526 243 528 245
rect 536 250 538 252
rect 536 243 538 245
rect 546 256 548 258
rect 546 249 548 251
rect 556 250 558 252
rect 556 243 558 245
rect 576 250 578 252
rect 576 243 578 245
rect 586 256 588 258
rect 586 249 588 251
rect 596 250 598 252
rect 596 243 598 245
rect 627 250 629 252
rect 627 243 629 245
rect 637 258 639 260
rect 637 251 639 253
rect 649 250 651 252
rect 649 243 651 245
rect 672 262 674 264
rect 684 243 686 245
rect 50 219 52 221
rect 71 225 73 227
rect 71 218 73 220
rect 81 217 83 219
rect 81 210 83 212
rect 93 225 95 227
rect 93 218 95 220
rect 128 225 130 227
rect 116 206 118 208
rect 172 225 174 227
rect 172 218 174 220
rect 182 217 184 219
rect 182 210 184 212
rect 194 225 196 227
rect 194 218 196 220
rect 229 225 231 227
rect 217 206 219 208
rect 274 225 276 227
rect 274 218 276 220
rect 284 217 286 219
rect 284 210 286 212
rect 296 225 298 227
rect 296 218 298 220
rect 331 225 333 227
rect 319 206 321 208
rect 394 219 396 221
rect 427 225 429 227
rect 427 218 429 220
rect 437 217 439 219
rect 437 210 439 212
rect 449 225 451 227
rect 449 218 451 220
rect 484 225 486 227
rect 472 206 474 208
rect 528 225 530 227
rect 528 218 530 220
rect 538 217 540 219
rect 538 210 540 212
rect 550 225 552 227
rect 550 218 552 220
rect 585 225 587 227
rect 573 206 575 208
rect 627 225 629 227
rect 627 218 629 220
rect 637 217 639 219
rect 637 210 639 212
rect 649 225 651 227
rect 649 218 651 220
rect 684 225 686 227
rect 672 206 674 208
rect 32 106 34 108
rect 32 99 34 101
rect 42 114 44 116
rect 42 107 44 109
rect 54 106 56 108
rect 54 99 56 101
rect 77 118 79 120
rect 89 99 91 101
rect 140 105 142 107
rect 173 106 175 108
rect 173 99 175 101
rect 183 114 185 116
rect 183 107 185 109
rect 195 106 197 108
rect 195 99 197 101
rect 218 118 220 120
rect 230 99 232 101
rect 286 118 288 120
rect 274 99 276 101
rect 309 106 311 108
rect 309 99 311 101
rect 321 114 323 116
rect 321 107 323 109
rect 331 106 333 108
rect 331 99 333 101
rect 394 105 396 107
rect 427 106 429 108
rect 427 99 429 101
rect 437 114 439 116
rect 437 107 439 109
rect 449 106 451 108
rect 449 99 451 101
rect 472 118 474 120
rect 484 99 486 101
rect 528 106 530 108
rect 528 99 530 101
rect 538 114 540 116
rect 538 107 540 109
rect 550 106 552 108
rect 550 99 552 101
rect 573 118 575 120
rect 585 99 587 101
rect 627 106 629 108
rect 627 99 629 101
rect 637 114 639 116
rect 637 107 639 109
rect 649 106 651 108
rect 649 99 651 101
rect 672 118 674 120
rect 684 99 686 101
rect 50 75 52 77
rect 71 81 73 83
rect 71 74 73 76
rect 81 73 83 75
rect 81 66 83 68
rect 93 81 95 83
rect 93 74 95 76
rect 128 81 130 83
rect 116 62 118 64
rect 172 81 174 83
rect 172 74 174 76
rect 182 73 184 75
rect 182 66 184 68
rect 194 81 196 83
rect 194 74 196 76
rect 229 81 231 83
rect 217 62 219 64
rect 273 81 275 83
rect 273 74 275 76
rect 283 73 285 75
rect 283 66 285 68
rect 295 81 297 83
rect 295 74 297 76
rect 330 81 332 83
rect 318 62 320 64
rect 393 75 395 77
rect 426 81 428 83
rect 426 74 428 76
rect 436 73 438 75
rect 436 66 438 68
rect 448 81 450 83
rect 448 74 450 76
rect 483 81 485 83
rect 471 62 473 64
rect 527 81 529 83
rect 527 74 529 76
rect 537 73 539 75
rect 537 66 539 68
rect 549 81 551 83
rect 549 74 551 76
rect 584 81 586 83
rect 572 62 574 64
rect 626 81 628 83
rect 626 74 628 76
rect 636 73 638 75
rect 636 66 638 68
rect 648 81 650 83
rect 648 74 650 76
rect 683 81 685 83
rect 671 62 673 64
<< pdifct1 >>
rect 50 362 52 364
rect 50 355 52 357
rect 90 362 92 364
rect 90 355 92 357
rect 101 354 103 356
rect 101 347 103 349
rect 179 357 181 359
rect 179 350 181 352
rect 197 357 199 359
rect 197 350 199 352
rect 286 362 288 364
rect 275 354 277 356
rect 286 355 288 357
rect 275 347 277 349
rect 326 362 328 364
rect 326 355 328 357
rect 367 357 369 359
rect 367 350 369 352
rect 456 362 458 364
rect 445 354 447 356
rect 456 355 458 357
rect 445 347 447 349
rect 496 362 498 364
rect 496 355 498 357
rect 566 362 568 364
rect 566 355 568 357
rect 606 362 608 364
rect 606 355 608 357
rect 617 354 619 356
rect 617 347 619 349
rect 695 357 697 359
rect 695 350 697 352
rect 50 257 52 259
rect 50 250 52 252
rect 101 265 103 267
rect 90 257 92 259
rect 90 250 92 252
rect 179 262 181 264
rect 179 255 181 257
rect 197 262 199 264
rect 197 255 199 257
rect 275 265 277 267
rect 275 258 277 260
rect 286 257 288 259
rect 286 250 288 252
rect 326 257 328 259
rect 326 250 328 252
rect 367 262 369 264
rect 367 255 369 257
rect 445 265 447 267
rect 445 258 447 260
rect 456 257 458 259
rect 456 250 458 252
rect 496 257 498 259
rect 496 250 498 252
rect 566 257 568 259
rect 566 250 568 252
rect 617 265 619 267
rect 606 257 608 259
rect 617 258 619 260
rect 606 250 608 252
rect 695 262 697 264
rect 695 255 697 257
rect 20 219 22 221
rect 20 212 22 214
rect 31 228 33 230
rect 61 210 63 212
rect 61 203 63 205
rect 139 213 141 215
rect 139 206 141 208
rect 162 210 164 212
rect 162 203 164 205
rect 240 213 242 215
rect 240 206 242 208
rect 264 210 266 212
rect 264 203 266 205
rect 364 219 366 221
rect 342 213 344 215
rect 364 212 366 214
rect 342 206 344 208
rect 375 228 377 230
rect 417 210 419 212
rect 417 203 419 205
rect 495 213 497 215
rect 495 206 497 208
rect 518 210 520 212
rect 518 203 520 205
rect 596 213 598 215
rect 596 206 598 208
rect 617 210 619 212
rect 617 203 619 205
rect 695 213 697 215
rect 695 206 697 208
rect 22 121 24 123
rect 22 114 24 116
rect 100 118 102 120
rect 100 111 102 113
rect 110 112 112 114
rect 110 105 112 107
rect 121 96 123 98
rect 163 121 165 123
rect 163 114 165 116
rect 241 118 243 120
rect 241 111 243 113
rect 263 118 265 120
rect 263 111 265 113
rect 341 121 343 123
rect 341 114 343 116
rect 364 112 366 114
rect 364 105 366 107
rect 375 96 377 98
rect 417 121 419 123
rect 417 114 419 116
rect 495 118 497 120
rect 495 111 497 113
rect 518 121 520 123
rect 518 114 520 116
rect 596 118 598 120
rect 596 111 598 113
rect 617 121 619 123
rect 617 114 619 116
rect 695 118 697 120
rect 695 111 697 113
rect 20 75 22 77
rect 20 68 22 70
rect 31 84 33 86
rect 61 66 63 68
rect 61 59 63 61
rect 139 69 141 71
rect 139 62 141 64
rect 162 66 164 68
rect 162 59 164 61
rect 240 69 242 71
rect 240 62 242 64
rect 263 66 265 68
rect 263 59 265 61
rect 363 75 365 77
rect 341 69 343 71
rect 363 68 365 70
rect 341 62 343 64
rect 374 84 376 86
rect 416 66 418 68
rect 416 59 418 61
rect 494 69 496 71
rect 494 62 496 64
rect 517 66 519 68
rect 517 59 519 61
rect 595 69 597 71
rect 595 62 597 64
rect 616 66 618 68
rect 616 59 618 61
rect 694 69 696 71
rect 694 62 696 64
<< alu0 >>
rect 18 369 20 371
rect 22 369 24 371
rect 18 364 24 369
rect 38 369 40 371
rect 42 369 44 371
rect 18 362 20 364
rect 22 362 24 364
rect 18 361 24 362
rect 28 365 34 366
rect 28 363 30 365
rect 32 363 34 365
rect 28 358 34 363
rect 38 364 44 369
rect 58 369 60 371
rect 62 369 64 371
rect 38 362 40 364
rect 42 362 44 364
rect 38 361 44 362
rect 28 356 30 358
rect 32 357 34 358
rect 58 364 64 369
rect 78 369 80 371
rect 82 369 84 371
rect 58 362 60 364
rect 62 362 64 364
rect 58 361 64 362
rect 68 365 74 366
rect 68 363 70 365
rect 72 363 74 365
rect 68 358 74 363
rect 78 364 84 369
rect 109 369 111 371
rect 113 369 115 371
rect 78 362 80 364
rect 82 362 84 364
rect 78 361 84 362
rect 32 356 42 357
rect 28 353 42 356
rect 38 349 42 353
rect 38 345 46 349
rect 42 340 46 345
rect 42 338 43 340
rect 45 338 46 340
rect 42 333 46 338
rect 34 329 46 333
rect 34 325 38 329
rect 49 326 50 333
rect 68 356 70 358
rect 72 357 74 358
rect 109 364 115 369
rect 131 369 133 371
rect 135 369 137 371
rect 109 362 111 364
rect 113 362 115 364
rect 109 361 115 362
rect 120 363 124 365
rect 120 361 121 363
rect 123 361 124 363
rect 131 364 137 369
rect 166 369 168 371
rect 170 369 172 371
rect 166 368 172 369
rect 206 369 208 371
rect 210 369 212 371
rect 206 368 212 369
rect 241 369 243 371
rect 245 369 247 371
rect 131 362 133 364
rect 135 362 137 364
rect 131 361 137 362
rect 72 356 82 357
rect 68 353 82 356
rect 78 349 82 353
rect 78 345 86 349
rect 82 340 86 345
rect 82 338 83 340
rect 85 338 86 340
rect 82 333 86 338
rect 74 329 86 333
rect 18 324 38 325
rect 18 322 20 324
rect 22 322 38 324
rect 18 321 38 322
rect 74 325 78 329
rect 89 326 90 333
rect 58 324 78 325
rect 58 322 60 324
rect 62 322 78 324
rect 58 321 78 322
rect 120 357 124 361
rect 143 357 167 361
rect 107 356 147 357
rect 107 354 121 356
rect 123 354 147 356
rect 107 353 147 354
rect 107 342 111 353
rect 155 352 159 354
rect 163 353 169 357
rect 155 350 156 352
rect 158 350 159 352
rect 155 349 159 350
rect 155 345 162 349
rect 105 340 111 342
rect 105 338 106 340
rect 108 338 111 340
rect 105 336 111 338
rect 115 340 119 345
rect 115 338 116 340
rect 118 338 119 340
rect 115 336 119 338
rect 107 333 111 336
rect 107 329 127 333
rect 123 325 127 329
rect 158 334 162 345
rect 165 343 169 353
rect 165 341 166 343
rect 168 341 169 343
rect 165 339 169 341
rect 158 333 176 334
rect 138 331 142 333
rect 158 332 172 333
rect 138 329 139 331
rect 141 329 142 331
rect 123 324 133 325
rect 123 322 129 324
rect 131 322 133 324
rect 123 321 133 322
rect 138 324 142 329
rect 147 331 172 332
rect 174 331 176 333
rect 147 329 149 331
rect 151 330 176 331
rect 151 329 162 330
rect 147 328 162 329
rect 138 322 139 324
rect 141 323 163 324
rect 141 322 159 323
rect 138 321 159 322
rect 161 321 163 323
rect 138 320 163 321
rect 168 320 172 322
rect 241 364 247 369
rect 263 369 265 371
rect 267 369 269 371
rect 241 362 243 364
rect 245 362 247 364
rect 241 361 247 362
rect 254 363 258 365
rect 254 361 255 363
rect 257 361 258 363
rect 263 364 269 369
rect 294 369 296 371
rect 298 369 300 371
rect 263 362 265 364
rect 267 362 269 364
rect 263 361 269 362
rect 211 357 235 361
rect 254 357 258 361
rect 209 353 215 357
rect 231 356 271 357
rect 231 354 255 356
rect 257 354 271 356
rect 209 343 213 353
rect 219 352 223 354
rect 231 353 271 354
rect 219 350 220 352
rect 222 350 223 352
rect 219 349 223 350
rect 209 341 210 343
rect 212 341 213 343
rect 209 339 213 341
rect 216 345 223 349
rect 216 334 220 345
rect 259 340 263 345
rect 259 338 260 340
rect 262 338 263 340
rect 202 333 220 334
rect 202 331 204 333
rect 206 332 220 333
rect 206 331 231 332
rect 202 330 227 331
rect 216 329 227 330
rect 229 329 231 331
rect 216 328 231 329
rect 236 331 240 333
rect 236 329 237 331
rect 239 329 240 331
rect 236 324 240 329
rect 259 336 263 338
rect 267 342 271 353
rect 267 340 273 342
rect 267 338 270 340
rect 272 338 273 340
rect 267 336 273 338
rect 267 333 271 336
rect 251 329 271 333
rect 251 325 255 329
rect 215 323 237 324
rect 206 320 210 322
rect 215 321 217 323
rect 219 322 237 323
rect 239 322 240 324
rect 219 321 240 322
rect 245 324 255 325
rect 245 322 247 324
rect 249 322 255 324
rect 245 321 255 322
rect 294 364 300 369
rect 314 369 316 371
rect 318 369 320 371
rect 294 362 296 364
rect 298 362 300 364
rect 294 361 300 362
rect 304 365 310 366
rect 304 363 306 365
rect 308 363 310 365
rect 304 358 310 363
rect 314 364 320 369
rect 334 369 336 371
rect 338 369 340 371
rect 314 362 316 364
rect 318 362 320 364
rect 314 361 320 362
rect 304 357 306 358
rect 296 356 306 357
rect 308 356 310 358
rect 296 353 310 356
rect 296 349 300 353
rect 292 345 300 349
rect 334 364 340 369
rect 354 369 356 371
rect 358 369 360 371
rect 334 362 336 364
rect 338 362 340 364
rect 334 361 340 362
rect 344 365 350 366
rect 344 363 346 365
rect 348 363 350 365
rect 344 358 350 363
rect 354 364 360 369
rect 376 369 378 371
rect 380 369 382 371
rect 376 368 382 369
rect 411 369 413 371
rect 415 369 417 371
rect 354 362 356 364
rect 358 362 360 364
rect 354 361 360 362
rect 411 364 417 369
rect 433 369 435 371
rect 437 369 439 371
rect 411 362 413 364
rect 415 362 417 364
rect 411 361 417 362
rect 424 363 428 365
rect 424 361 425 363
rect 427 361 428 363
rect 433 364 439 369
rect 464 369 466 371
rect 468 369 470 371
rect 433 362 435 364
rect 437 362 439 364
rect 433 361 439 362
rect 344 357 346 358
rect 336 356 346 357
rect 348 356 350 358
rect 336 353 350 356
rect 292 340 296 345
rect 292 338 293 340
rect 295 338 296 340
rect 292 333 296 338
rect 288 326 289 333
rect 292 329 304 333
rect 300 325 304 329
rect 336 349 340 353
rect 332 345 340 349
rect 381 357 405 361
rect 424 357 428 361
rect 379 353 385 357
rect 401 356 441 357
rect 401 354 425 356
rect 427 354 441 356
rect 332 340 336 345
rect 332 338 333 340
rect 335 338 336 340
rect 332 333 336 338
rect 328 326 329 333
rect 332 329 344 333
rect 300 324 320 325
rect 300 322 316 324
rect 318 322 320 324
rect 300 321 320 322
rect 340 325 344 329
rect 379 343 383 353
rect 389 352 393 354
rect 401 353 441 354
rect 389 350 390 352
rect 392 350 393 352
rect 389 349 393 350
rect 379 341 380 343
rect 382 341 383 343
rect 379 339 383 341
rect 386 345 393 349
rect 386 334 390 345
rect 429 340 433 345
rect 429 338 430 340
rect 432 338 433 340
rect 372 333 390 334
rect 372 331 374 333
rect 376 332 390 333
rect 376 331 401 332
rect 372 330 397 331
rect 386 329 397 330
rect 399 329 401 331
rect 386 328 401 329
rect 406 331 410 333
rect 406 329 407 331
rect 409 329 410 331
rect 340 324 360 325
rect 340 322 356 324
rect 358 322 360 324
rect 340 321 360 322
rect 406 324 410 329
rect 429 336 433 338
rect 437 342 441 353
rect 437 340 443 342
rect 437 338 440 340
rect 442 338 443 340
rect 437 336 443 338
rect 437 333 441 336
rect 421 329 441 333
rect 421 325 425 329
rect 385 323 407 324
rect 215 320 240 321
rect 376 320 380 322
rect 385 321 387 323
rect 389 322 407 323
rect 409 322 410 324
rect 389 321 410 322
rect 415 324 425 325
rect 415 322 417 324
rect 419 322 425 324
rect 415 321 425 322
rect 464 364 470 369
rect 484 369 486 371
rect 488 369 490 371
rect 464 362 466 364
rect 468 362 470 364
rect 464 361 470 362
rect 474 365 480 366
rect 474 363 476 365
rect 478 363 480 365
rect 474 358 480 363
rect 484 364 490 369
rect 504 369 506 371
rect 508 369 510 371
rect 484 362 486 364
rect 488 362 490 364
rect 484 361 490 362
rect 474 357 476 358
rect 466 356 476 357
rect 478 356 480 358
rect 466 353 480 356
rect 466 349 470 353
rect 462 345 470 349
rect 504 364 510 369
rect 524 369 526 371
rect 528 369 530 371
rect 504 362 506 364
rect 508 362 510 364
rect 504 361 510 362
rect 514 365 520 366
rect 514 363 516 365
rect 518 363 520 365
rect 514 358 520 363
rect 524 364 530 369
rect 524 362 526 364
rect 528 362 530 364
rect 524 361 530 362
rect 534 369 536 371
rect 538 369 540 371
rect 534 364 540 369
rect 554 369 556 371
rect 558 369 560 371
rect 534 362 536 364
rect 538 362 540 364
rect 534 361 540 362
rect 544 365 550 366
rect 544 363 546 365
rect 548 363 550 365
rect 544 358 550 363
rect 554 364 560 369
rect 574 369 576 371
rect 578 369 580 371
rect 554 362 556 364
rect 558 362 560 364
rect 554 361 560 362
rect 514 357 516 358
rect 506 356 516 357
rect 518 356 520 358
rect 506 353 520 356
rect 462 340 466 345
rect 462 338 463 340
rect 465 338 466 340
rect 462 333 466 338
rect 458 326 459 333
rect 462 329 474 333
rect 470 325 474 329
rect 506 349 510 353
rect 502 345 510 349
rect 544 356 546 358
rect 548 357 550 358
rect 574 364 580 369
rect 594 369 596 371
rect 598 369 600 371
rect 574 362 576 364
rect 578 362 580 364
rect 574 361 580 362
rect 584 365 590 366
rect 584 363 586 365
rect 588 363 590 365
rect 584 358 590 363
rect 594 364 600 369
rect 625 369 627 371
rect 629 369 631 371
rect 594 362 596 364
rect 598 362 600 364
rect 594 361 600 362
rect 548 356 558 357
rect 544 353 558 356
rect 554 349 558 353
rect 554 345 562 349
rect 502 340 506 345
rect 502 338 503 340
rect 505 338 506 340
rect 502 333 506 338
rect 498 326 499 333
rect 502 329 514 333
rect 470 324 490 325
rect 470 322 486 324
rect 488 322 490 324
rect 470 321 490 322
rect 510 325 514 329
rect 558 340 562 345
rect 558 338 559 340
rect 561 338 562 340
rect 558 333 562 338
rect 550 329 562 333
rect 550 325 554 329
rect 565 326 566 333
rect 584 356 586 358
rect 588 357 590 358
rect 625 364 631 369
rect 647 369 649 371
rect 651 369 653 371
rect 625 362 627 364
rect 629 362 631 364
rect 625 361 631 362
rect 636 363 640 365
rect 636 361 637 363
rect 639 361 640 363
rect 647 364 653 369
rect 682 369 684 371
rect 686 369 688 371
rect 682 368 688 369
rect 647 362 649 364
rect 651 362 653 364
rect 647 361 653 362
rect 588 356 598 357
rect 584 353 598 356
rect 594 349 598 353
rect 594 345 602 349
rect 598 340 602 345
rect 598 338 599 340
rect 601 338 602 340
rect 598 333 602 338
rect 590 329 602 333
rect 510 324 530 325
rect 510 322 526 324
rect 528 322 530 324
rect 510 321 530 322
rect 534 324 554 325
rect 534 322 536 324
rect 538 322 554 324
rect 534 321 554 322
rect 590 325 594 329
rect 605 326 606 333
rect 574 324 594 325
rect 574 322 576 324
rect 578 322 594 324
rect 574 321 594 322
rect 636 357 640 361
rect 659 357 683 361
rect 623 356 663 357
rect 623 354 637 356
rect 639 354 663 356
rect 623 353 663 354
rect 623 342 627 353
rect 671 352 675 354
rect 679 353 685 357
rect 671 350 672 352
rect 674 350 675 352
rect 671 349 675 350
rect 671 345 678 349
rect 621 340 627 342
rect 621 338 622 340
rect 624 338 627 340
rect 621 336 627 338
rect 631 340 635 345
rect 631 338 632 340
rect 634 338 635 340
rect 631 336 635 338
rect 623 333 627 336
rect 623 329 643 333
rect 639 325 643 329
rect 674 334 678 345
rect 681 343 685 353
rect 681 341 682 343
rect 684 341 685 343
rect 681 339 685 341
rect 674 333 692 334
rect 654 331 658 333
rect 674 332 688 333
rect 654 329 655 331
rect 657 329 658 331
rect 639 324 649 325
rect 639 322 645 324
rect 647 322 649 324
rect 639 321 649 322
rect 654 324 658 329
rect 663 331 688 332
rect 690 331 692 333
rect 663 329 665 331
rect 667 330 692 331
rect 667 329 678 330
rect 663 328 678 329
rect 654 322 655 324
rect 657 323 679 324
rect 657 322 675 323
rect 654 321 675 322
rect 677 321 679 323
rect 385 320 410 321
rect 654 320 679 321
rect 684 320 688 322
rect 168 318 169 320
rect 171 318 172 320
rect 110 317 116 318
rect 110 315 112 317
rect 114 315 116 317
rect 168 315 172 318
rect 206 318 207 320
rect 209 318 210 320
rect 376 318 377 320
rect 379 318 380 320
rect 684 318 685 320
rect 687 318 688 320
rect 206 315 210 318
rect 262 317 268 318
rect 262 315 264 317
rect 266 315 268 317
rect 376 315 380 318
rect 432 317 438 318
rect 432 315 434 317
rect 436 315 438 317
rect 626 317 632 318
rect 626 315 628 317
rect 630 315 632 317
rect 684 315 688 318
rect 110 297 112 299
rect 114 297 116 299
rect 110 296 116 297
rect 168 296 172 299
rect 168 294 169 296
rect 171 294 172 296
rect 206 296 210 299
rect 262 297 264 299
rect 266 297 268 299
rect 262 296 268 297
rect 376 296 380 299
rect 432 297 434 299
rect 436 297 438 299
rect 432 296 438 297
rect 626 297 628 299
rect 630 297 632 299
rect 626 296 632 297
rect 684 296 688 299
rect 206 294 207 296
rect 209 294 210 296
rect 376 294 377 296
rect 379 294 380 296
rect 684 294 685 296
rect 687 294 688 296
rect 138 293 163 294
rect 18 292 38 293
rect 18 290 20 292
rect 22 290 38 292
rect 18 289 38 290
rect 34 285 38 289
rect 58 292 78 293
rect 58 290 60 292
rect 62 290 78 292
rect 58 289 78 290
rect 34 281 46 285
rect 49 281 50 288
rect 42 276 46 281
rect 42 274 43 276
rect 45 274 46 276
rect 42 269 46 274
rect 38 265 46 269
rect 38 261 42 265
rect 74 285 78 289
rect 74 281 86 285
rect 89 281 90 288
rect 82 276 86 281
rect 82 274 83 276
rect 85 274 86 276
rect 82 269 86 274
rect 28 258 42 261
rect 28 256 30 258
rect 32 257 42 258
rect 32 256 34 257
rect 18 252 24 253
rect 18 250 20 252
rect 22 250 24 252
rect 18 245 24 250
rect 28 251 34 256
rect 28 249 30 251
rect 32 249 34 251
rect 28 248 34 249
rect 38 252 44 253
rect 38 250 40 252
rect 42 250 44 252
rect 18 243 20 245
rect 22 243 24 245
rect 38 245 44 250
rect 78 265 86 269
rect 78 261 82 265
rect 68 258 82 261
rect 68 256 70 258
rect 72 257 82 258
rect 72 256 74 257
rect 58 252 64 253
rect 58 250 60 252
rect 62 250 64 252
rect 38 243 40 245
rect 42 243 44 245
rect 58 245 64 250
rect 68 251 74 256
rect 68 249 70 251
rect 72 249 74 251
rect 68 248 74 249
rect 78 252 84 253
rect 78 250 80 252
rect 82 250 84 252
rect 58 243 60 245
rect 62 243 64 245
rect 78 245 84 250
rect 123 292 133 293
rect 123 290 129 292
rect 131 290 133 292
rect 123 289 133 290
rect 138 292 159 293
rect 138 290 139 292
rect 141 291 159 292
rect 161 291 163 293
rect 168 292 172 294
rect 141 290 163 291
rect 123 285 127 289
rect 107 281 127 285
rect 107 278 111 281
rect 105 276 111 278
rect 105 274 106 276
rect 108 274 111 276
rect 105 272 111 274
rect 100 260 104 261
rect 100 258 101 260
rect 103 258 104 260
rect 100 257 104 258
rect 107 261 111 272
rect 115 276 119 278
rect 138 285 142 290
rect 138 283 139 285
rect 141 283 142 285
rect 138 281 142 283
rect 147 285 162 286
rect 147 283 149 285
rect 151 284 162 285
rect 151 283 176 284
rect 147 282 172 283
rect 158 281 172 282
rect 174 281 176 283
rect 158 280 176 281
rect 115 274 116 276
rect 118 274 119 276
rect 115 269 119 274
rect 158 269 162 280
rect 155 265 162 269
rect 165 273 169 275
rect 165 271 166 273
rect 168 271 169 273
rect 155 264 159 265
rect 155 262 156 264
rect 158 262 159 264
rect 107 260 147 261
rect 155 260 159 262
rect 165 261 169 271
rect 107 258 121 260
rect 123 258 147 260
rect 107 257 147 258
rect 163 257 169 261
rect 120 253 124 257
rect 143 253 167 257
rect 109 252 115 253
rect 109 250 111 252
rect 113 250 115 252
rect 78 243 80 245
rect 82 243 84 245
rect 109 245 115 250
rect 120 251 121 253
rect 123 251 124 253
rect 120 249 124 251
rect 131 252 137 253
rect 131 250 133 252
rect 135 250 137 252
rect 109 243 111 245
rect 113 243 115 245
rect 131 245 137 250
rect 206 292 210 294
rect 215 293 240 294
rect 215 291 217 293
rect 219 292 240 293
rect 219 291 237 292
rect 215 290 237 291
rect 239 290 240 292
rect 216 285 231 286
rect 216 284 227 285
rect 202 283 227 284
rect 229 283 231 285
rect 202 281 204 283
rect 206 282 231 283
rect 236 285 240 290
rect 245 292 255 293
rect 245 290 247 292
rect 249 290 255 292
rect 245 289 255 290
rect 236 283 237 285
rect 239 283 240 285
rect 206 281 220 282
rect 236 281 240 283
rect 202 280 220 281
rect 209 273 213 275
rect 209 271 210 273
rect 212 271 213 273
rect 209 261 213 271
rect 216 269 220 280
rect 251 285 255 289
rect 251 281 271 285
rect 267 278 271 281
rect 259 276 263 278
rect 259 274 260 276
rect 262 274 263 276
rect 259 269 263 274
rect 267 276 273 278
rect 267 274 270 276
rect 272 274 273 276
rect 267 272 273 274
rect 216 265 223 269
rect 219 264 223 265
rect 219 262 220 264
rect 222 262 223 264
rect 209 257 215 261
rect 219 260 223 262
rect 267 261 271 272
rect 231 260 271 261
rect 231 258 255 260
rect 257 258 271 260
rect 231 257 271 258
rect 211 253 235 257
rect 254 253 258 257
rect 300 292 320 293
rect 300 290 316 292
rect 318 290 320 292
rect 300 289 320 290
rect 288 281 289 288
rect 300 285 304 289
rect 340 292 360 293
rect 340 290 356 292
rect 358 290 360 292
rect 340 289 360 290
rect 376 292 380 294
rect 385 293 410 294
rect 654 293 679 294
rect 385 291 387 293
rect 389 292 410 293
rect 389 291 407 292
rect 385 290 407 291
rect 409 290 410 292
rect 292 281 304 285
rect 292 276 296 281
rect 292 274 293 276
rect 295 274 296 276
rect 292 269 296 274
rect 292 265 300 269
rect 296 261 300 265
rect 296 258 310 261
rect 296 257 306 258
rect 241 252 247 253
rect 241 250 243 252
rect 245 250 247 252
rect 131 243 133 245
rect 135 243 137 245
rect 166 245 172 246
rect 166 243 168 245
rect 170 243 172 245
rect 206 245 212 246
rect 206 243 208 245
rect 210 243 212 245
rect 241 245 247 250
rect 254 251 255 253
rect 257 251 258 253
rect 254 249 258 251
rect 263 252 269 253
rect 263 250 265 252
rect 267 250 269 252
rect 241 243 243 245
rect 245 243 247 245
rect 263 245 269 250
rect 304 256 306 257
rect 308 256 310 258
rect 328 281 329 288
rect 340 285 344 289
rect 332 281 344 285
rect 332 276 336 281
rect 332 274 333 276
rect 335 274 336 276
rect 332 269 336 274
rect 332 265 340 269
rect 336 261 340 265
rect 336 258 350 261
rect 336 257 346 258
rect 294 252 300 253
rect 294 250 296 252
rect 298 250 300 252
rect 263 243 265 245
rect 267 243 269 245
rect 294 245 300 250
rect 304 251 310 256
rect 344 256 346 257
rect 348 256 350 258
rect 386 285 401 286
rect 386 284 397 285
rect 372 283 397 284
rect 399 283 401 285
rect 372 281 374 283
rect 376 282 401 283
rect 406 285 410 290
rect 415 292 425 293
rect 415 290 417 292
rect 419 290 425 292
rect 415 289 425 290
rect 406 283 407 285
rect 409 283 410 285
rect 376 281 390 282
rect 406 281 410 283
rect 372 280 390 281
rect 379 273 383 275
rect 379 271 380 273
rect 382 271 383 273
rect 379 261 383 271
rect 386 269 390 280
rect 421 285 425 289
rect 421 281 441 285
rect 437 278 441 281
rect 429 276 433 278
rect 429 274 430 276
rect 432 274 433 276
rect 429 269 433 274
rect 437 276 443 278
rect 437 274 440 276
rect 442 274 443 276
rect 437 272 443 274
rect 386 265 393 269
rect 389 264 393 265
rect 389 262 390 264
rect 392 262 393 264
rect 379 257 385 261
rect 389 260 393 262
rect 437 261 441 272
rect 401 260 441 261
rect 401 258 425 260
rect 427 258 441 260
rect 401 257 441 258
rect 304 249 306 251
rect 308 249 310 251
rect 304 248 310 249
rect 314 252 320 253
rect 314 250 316 252
rect 318 250 320 252
rect 294 243 296 245
rect 298 243 300 245
rect 314 245 320 250
rect 334 252 340 253
rect 334 250 336 252
rect 338 250 340 252
rect 314 243 316 245
rect 318 243 320 245
rect 334 245 340 250
rect 344 251 350 256
rect 381 253 405 257
rect 424 253 428 257
rect 470 292 490 293
rect 470 290 486 292
rect 488 290 490 292
rect 470 289 490 290
rect 458 281 459 288
rect 470 285 474 289
rect 510 292 530 293
rect 510 290 526 292
rect 528 290 530 292
rect 510 289 530 290
rect 534 292 554 293
rect 534 290 536 292
rect 538 290 554 292
rect 534 289 554 290
rect 462 281 474 285
rect 462 276 466 281
rect 462 274 463 276
rect 465 274 466 276
rect 462 269 466 274
rect 498 281 499 288
rect 510 285 514 289
rect 502 281 514 285
rect 462 265 470 269
rect 466 261 470 265
rect 466 258 480 261
rect 466 257 476 258
rect 344 249 346 251
rect 348 249 350 251
rect 344 248 350 249
rect 354 252 360 253
rect 354 250 356 252
rect 358 250 360 252
rect 334 243 336 245
rect 338 243 340 245
rect 354 245 360 250
rect 411 252 417 253
rect 411 250 413 252
rect 415 250 417 252
rect 354 243 356 245
rect 358 243 360 245
rect 376 245 382 246
rect 376 243 378 245
rect 380 243 382 245
rect 411 245 417 250
rect 424 251 425 253
rect 427 251 428 253
rect 424 249 428 251
rect 433 252 439 253
rect 433 250 435 252
rect 437 250 439 252
rect 411 243 413 245
rect 415 243 417 245
rect 433 245 439 250
rect 474 256 476 257
rect 478 256 480 258
rect 502 276 506 281
rect 502 274 503 276
rect 505 274 506 276
rect 502 269 506 274
rect 550 285 554 289
rect 574 292 594 293
rect 574 290 576 292
rect 578 290 594 292
rect 574 289 594 290
rect 550 281 562 285
rect 565 281 566 288
rect 558 276 562 281
rect 558 274 559 276
rect 561 274 562 276
rect 558 269 562 274
rect 502 265 510 269
rect 506 261 510 265
rect 506 258 520 261
rect 506 257 516 258
rect 464 252 470 253
rect 464 250 466 252
rect 468 250 470 252
rect 433 243 435 245
rect 437 243 439 245
rect 464 245 470 250
rect 474 251 480 256
rect 474 249 476 251
rect 478 249 480 251
rect 474 248 480 249
rect 484 252 490 253
rect 484 250 486 252
rect 488 250 490 252
rect 464 243 466 245
rect 468 243 470 245
rect 484 245 490 250
rect 514 256 516 257
rect 518 256 520 258
rect 554 265 562 269
rect 554 261 558 265
rect 590 285 594 289
rect 590 281 602 285
rect 605 281 606 288
rect 598 276 602 281
rect 598 274 599 276
rect 601 274 602 276
rect 598 269 602 274
rect 544 258 558 261
rect 544 256 546 258
rect 548 257 558 258
rect 548 256 550 257
rect 504 252 510 253
rect 504 250 506 252
rect 508 250 510 252
rect 484 243 486 245
rect 488 243 490 245
rect 504 245 510 250
rect 514 251 520 256
rect 514 249 516 251
rect 518 249 520 251
rect 514 248 520 249
rect 524 252 530 253
rect 524 250 526 252
rect 528 250 530 252
rect 504 243 506 245
rect 508 243 510 245
rect 524 245 530 250
rect 524 243 526 245
rect 528 243 530 245
rect 534 252 540 253
rect 534 250 536 252
rect 538 250 540 252
rect 534 245 540 250
rect 544 251 550 256
rect 544 249 546 251
rect 548 249 550 251
rect 544 248 550 249
rect 554 252 560 253
rect 554 250 556 252
rect 558 250 560 252
rect 534 243 536 245
rect 538 243 540 245
rect 554 245 560 250
rect 594 265 602 269
rect 594 261 598 265
rect 584 258 598 261
rect 584 256 586 258
rect 588 257 598 258
rect 588 256 590 257
rect 574 252 580 253
rect 574 250 576 252
rect 578 250 580 252
rect 554 243 556 245
rect 558 243 560 245
rect 574 245 580 250
rect 584 251 590 256
rect 584 249 586 251
rect 588 249 590 251
rect 584 248 590 249
rect 594 252 600 253
rect 594 250 596 252
rect 598 250 600 252
rect 574 243 576 245
rect 578 243 580 245
rect 594 245 600 250
rect 639 292 649 293
rect 639 290 645 292
rect 647 290 649 292
rect 639 289 649 290
rect 654 292 675 293
rect 654 290 655 292
rect 657 291 675 292
rect 677 291 679 293
rect 684 292 688 294
rect 657 290 679 291
rect 639 285 643 289
rect 623 281 643 285
rect 623 278 627 281
rect 621 276 627 278
rect 621 274 622 276
rect 624 274 627 276
rect 621 272 627 274
rect 623 261 627 272
rect 631 276 635 278
rect 654 285 658 290
rect 654 283 655 285
rect 657 283 658 285
rect 654 281 658 283
rect 663 285 678 286
rect 663 283 665 285
rect 667 284 678 285
rect 667 283 692 284
rect 663 282 688 283
rect 674 281 688 282
rect 690 281 692 283
rect 674 280 692 281
rect 631 274 632 276
rect 634 274 635 276
rect 631 269 635 274
rect 674 269 678 280
rect 671 265 678 269
rect 681 273 685 275
rect 681 271 682 273
rect 684 271 685 273
rect 671 264 675 265
rect 671 262 672 264
rect 674 262 675 264
rect 623 260 663 261
rect 671 260 675 262
rect 681 261 685 271
rect 623 258 637 260
rect 639 258 663 260
rect 623 257 663 258
rect 679 257 685 261
rect 636 253 640 257
rect 659 253 683 257
rect 625 252 631 253
rect 625 250 627 252
rect 629 250 631 252
rect 594 243 596 245
rect 598 243 600 245
rect 625 245 631 250
rect 636 251 637 253
rect 639 251 640 253
rect 636 249 640 251
rect 647 252 653 253
rect 647 250 649 252
rect 651 250 653 252
rect 625 243 627 245
rect 629 243 631 245
rect 647 245 653 250
rect 647 243 649 245
rect 651 243 653 245
rect 682 245 688 246
rect 682 243 684 245
rect 686 243 688 245
rect 69 225 71 227
rect 73 225 75 227
rect 34 221 54 222
rect 34 219 50 221
rect 52 219 54 221
rect 34 218 54 219
rect 69 220 75 225
rect 91 225 93 227
rect 95 225 97 227
rect 69 218 71 220
rect 73 218 75 220
rect 22 210 23 216
rect 34 213 38 218
rect 69 217 75 218
rect 80 219 84 221
rect 80 217 81 219
rect 83 217 84 219
rect 91 220 97 225
rect 126 225 128 227
rect 130 225 132 227
rect 126 224 132 225
rect 170 225 172 227
rect 174 225 176 227
rect 91 218 93 220
rect 95 218 97 220
rect 91 217 97 218
rect 170 220 176 225
rect 192 225 194 227
rect 196 225 198 227
rect 170 218 172 220
rect 174 218 176 220
rect 170 217 176 218
rect 181 219 185 221
rect 181 217 182 219
rect 184 217 185 219
rect 192 220 198 225
rect 227 225 229 227
rect 231 225 233 227
rect 227 224 233 225
rect 272 225 274 227
rect 276 225 278 227
rect 192 218 194 220
rect 196 218 198 220
rect 192 217 198 218
rect 272 220 278 225
rect 294 225 296 227
rect 298 225 300 227
rect 272 218 274 220
rect 276 218 278 220
rect 272 217 278 218
rect 283 219 287 221
rect 283 217 284 219
rect 286 217 287 219
rect 294 220 300 225
rect 329 225 331 227
rect 333 225 335 227
rect 329 224 335 225
rect 425 225 427 227
rect 429 225 431 227
rect 294 218 296 220
rect 298 218 300 220
rect 294 217 300 218
rect 26 209 38 213
rect 80 213 84 217
rect 103 213 127 217
rect 26 196 30 209
rect 26 194 27 196
rect 29 194 30 196
rect 26 188 30 194
rect 49 192 50 208
rect 67 212 107 213
rect 67 210 81 212
rect 83 210 107 212
rect 67 209 107 210
rect 26 184 43 188
rect 39 182 43 184
rect 28 180 34 181
rect 28 178 30 180
rect 32 178 34 180
rect 39 180 40 182
rect 42 180 43 182
rect 39 178 43 180
rect 48 182 54 183
rect 48 180 50 182
rect 52 180 54 182
rect 28 171 34 178
rect 48 171 54 180
rect 67 198 71 209
rect 115 208 119 210
rect 123 209 129 213
rect 115 206 116 208
rect 118 206 119 208
rect 115 205 119 206
rect 115 201 122 205
rect 65 196 71 198
rect 65 194 66 196
rect 68 194 71 196
rect 65 192 71 194
rect 75 196 79 201
rect 75 194 76 196
rect 78 194 79 196
rect 75 192 79 194
rect 67 189 71 192
rect 67 185 87 189
rect 83 181 87 185
rect 118 190 122 201
rect 125 199 129 209
rect 125 197 126 199
rect 128 197 129 199
rect 125 195 129 197
rect 118 189 136 190
rect 98 187 102 189
rect 118 188 132 189
rect 98 185 99 187
rect 101 185 102 187
rect 83 180 93 181
rect 83 178 89 180
rect 91 178 93 180
rect 83 177 93 178
rect 98 180 102 185
rect 107 187 132 188
rect 134 187 136 189
rect 107 185 109 187
rect 111 186 136 187
rect 111 185 122 186
rect 107 184 122 185
rect 98 178 99 180
rect 101 179 123 180
rect 101 178 119 179
rect 98 177 119 178
rect 121 177 123 179
rect 98 176 123 177
rect 128 176 132 178
rect 181 213 185 217
rect 204 213 228 217
rect 168 212 208 213
rect 168 210 182 212
rect 184 210 208 212
rect 168 209 208 210
rect 168 198 172 209
rect 216 208 220 210
rect 224 209 230 213
rect 216 206 217 208
rect 219 206 220 208
rect 216 205 220 206
rect 216 201 223 205
rect 166 196 172 198
rect 166 194 167 196
rect 169 194 172 196
rect 166 192 172 194
rect 176 196 180 201
rect 176 194 177 196
rect 179 194 180 196
rect 176 192 180 194
rect 168 189 172 192
rect 168 185 188 189
rect 184 181 188 185
rect 219 190 223 201
rect 226 199 230 209
rect 226 197 227 199
rect 229 197 230 199
rect 226 195 230 197
rect 219 189 237 190
rect 199 187 203 189
rect 219 188 233 189
rect 199 185 200 187
rect 202 185 203 187
rect 184 180 194 181
rect 184 178 190 180
rect 192 178 194 180
rect 184 177 194 178
rect 199 180 203 185
rect 208 187 233 188
rect 235 187 237 189
rect 208 185 210 187
rect 212 186 237 187
rect 212 185 223 186
rect 208 184 223 185
rect 199 178 200 180
rect 202 179 224 180
rect 202 178 220 179
rect 199 177 220 178
rect 222 177 224 179
rect 199 176 224 177
rect 229 176 233 178
rect 283 213 287 217
rect 306 213 330 217
rect 270 212 310 213
rect 270 210 284 212
rect 286 210 310 212
rect 270 209 310 210
rect 270 198 274 209
rect 318 208 322 210
rect 326 209 332 213
rect 318 206 319 208
rect 321 206 322 208
rect 318 205 322 206
rect 318 201 325 205
rect 268 196 274 198
rect 268 194 269 196
rect 271 194 274 196
rect 268 192 274 194
rect 278 196 282 201
rect 278 194 279 196
rect 281 194 282 196
rect 278 192 282 194
rect 270 189 274 192
rect 270 185 290 189
rect 286 181 290 185
rect 321 190 325 201
rect 328 199 332 209
rect 328 197 329 199
rect 331 197 332 199
rect 328 195 332 197
rect 321 189 339 190
rect 301 187 305 189
rect 321 188 335 189
rect 301 185 302 187
rect 304 185 305 187
rect 286 180 296 181
rect 286 178 292 180
rect 294 178 296 180
rect 286 177 296 178
rect 301 180 305 185
rect 310 187 335 188
rect 337 187 339 189
rect 310 185 312 187
rect 314 186 339 187
rect 314 185 325 186
rect 310 184 325 185
rect 301 178 302 180
rect 304 179 326 180
rect 304 178 322 179
rect 301 177 322 178
rect 324 177 326 179
rect 301 176 326 177
rect 331 176 335 178
rect 378 221 398 222
rect 378 219 394 221
rect 396 219 398 221
rect 378 218 398 219
rect 425 220 431 225
rect 447 225 449 227
rect 451 225 453 227
rect 425 218 427 220
rect 429 218 431 220
rect 366 210 367 216
rect 378 213 382 218
rect 425 217 431 218
rect 436 219 440 221
rect 436 217 437 219
rect 439 217 440 219
rect 447 220 453 225
rect 482 225 484 227
rect 486 225 488 227
rect 482 224 488 225
rect 526 225 528 227
rect 530 225 532 227
rect 447 218 449 220
rect 451 218 453 220
rect 447 217 453 218
rect 526 220 532 225
rect 548 225 550 227
rect 552 225 554 227
rect 526 218 528 220
rect 530 218 532 220
rect 526 217 532 218
rect 537 219 541 221
rect 537 217 538 219
rect 540 217 541 219
rect 548 220 554 225
rect 583 225 585 227
rect 587 225 589 227
rect 583 224 589 225
rect 625 225 627 227
rect 629 225 631 227
rect 548 218 550 220
rect 552 218 554 220
rect 548 217 554 218
rect 625 220 631 225
rect 647 225 649 227
rect 651 225 653 227
rect 625 218 627 220
rect 629 218 631 220
rect 625 217 631 218
rect 636 219 640 221
rect 636 217 637 219
rect 639 217 640 219
rect 647 220 653 225
rect 682 225 684 227
rect 686 225 688 227
rect 682 224 688 225
rect 647 218 649 220
rect 651 218 653 220
rect 647 217 653 218
rect 370 209 382 213
rect 436 213 440 217
rect 459 213 483 217
rect 370 196 374 209
rect 370 194 371 196
rect 373 194 374 196
rect 370 188 374 194
rect 393 192 394 208
rect 423 212 463 213
rect 423 210 437 212
rect 439 210 463 212
rect 423 209 463 210
rect 370 184 387 188
rect 383 182 387 184
rect 372 180 378 181
rect 372 178 374 180
rect 376 178 378 180
rect 383 180 384 182
rect 386 180 387 182
rect 383 178 387 180
rect 392 182 398 183
rect 392 180 394 182
rect 396 180 398 182
rect 128 174 129 176
rect 131 174 132 176
rect 229 174 230 176
rect 232 174 233 176
rect 331 174 332 176
rect 334 174 335 176
rect 70 173 76 174
rect 70 171 72 173
rect 74 171 76 173
rect 128 171 132 174
rect 171 173 177 174
rect 171 171 173 173
rect 175 171 177 173
rect 229 171 233 174
rect 273 173 279 174
rect 273 171 275 173
rect 277 171 279 173
rect 331 171 335 174
rect 372 171 378 178
rect 392 171 398 180
rect 423 198 427 209
rect 471 208 475 210
rect 479 209 485 213
rect 471 206 472 208
rect 474 206 475 208
rect 471 205 475 206
rect 471 201 478 205
rect 421 196 427 198
rect 421 194 422 196
rect 424 194 427 196
rect 421 192 427 194
rect 431 196 435 201
rect 431 194 432 196
rect 434 194 435 196
rect 431 192 435 194
rect 423 189 427 192
rect 423 185 443 189
rect 439 181 443 185
rect 474 190 478 201
rect 481 199 485 209
rect 481 197 482 199
rect 484 197 485 199
rect 481 195 485 197
rect 474 189 492 190
rect 454 187 458 189
rect 474 188 488 189
rect 454 185 455 187
rect 457 185 458 187
rect 439 180 449 181
rect 439 178 445 180
rect 447 178 449 180
rect 439 177 449 178
rect 454 180 458 185
rect 463 187 488 188
rect 490 187 492 189
rect 463 185 465 187
rect 467 186 492 187
rect 467 185 478 186
rect 463 184 478 185
rect 454 178 455 180
rect 457 179 479 180
rect 457 178 475 179
rect 454 177 475 178
rect 477 177 479 179
rect 454 176 479 177
rect 484 176 488 178
rect 537 213 541 217
rect 560 213 584 217
rect 524 212 564 213
rect 524 210 538 212
rect 540 210 564 212
rect 524 209 564 210
rect 524 198 528 209
rect 572 208 576 210
rect 580 209 586 213
rect 572 206 573 208
rect 575 206 576 208
rect 572 205 576 206
rect 572 201 579 205
rect 522 196 528 198
rect 522 194 523 196
rect 525 194 528 196
rect 522 192 528 194
rect 532 196 536 201
rect 532 194 533 196
rect 535 194 536 196
rect 532 192 536 194
rect 524 189 528 192
rect 524 185 544 189
rect 540 181 544 185
rect 575 190 579 201
rect 582 199 586 209
rect 582 197 583 199
rect 585 197 586 199
rect 582 195 586 197
rect 575 189 593 190
rect 555 187 559 189
rect 575 188 589 189
rect 555 185 556 187
rect 558 185 559 187
rect 540 180 550 181
rect 540 178 546 180
rect 548 178 550 180
rect 540 177 550 178
rect 555 180 559 185
rect 564 187 589 188
rect 591 187 593 189
rect 564 185 566 187
rect 568 186 593 187
rect 568 185 579 186
rect 564 184 579 185
rect 555 178 556 180
rect 558 179 580 180
rect 558 178 576 179
rect 555 177 576 178
rect 578 177 580 179
rect 555 176 580 177
rect 585 176 589 178
rect 636 213 640 217
rect 659 213 683 217
rect 623 212 663 213
rect 623 210 637 212
rect 639 210 663 212
rect 623 209 663 210
rect 623 198 627 209
rect 671 208 675 210
rect 679 209 685 213
rect 671 206 672 208
rect 674 206 675 208
rect 671 205 675 206
rect 671 201 678 205
rect 621 196 627 198
rect 621 194 622 196
rect 624 194 627 196
rect 621 192 627 194
rect 631 196 635 201
rect 631 194 632 196
rect 634 194 635 196
rect 631 192 635 194
rect 623 189 627 192
rect 623 185 643 189
rect 639 181 643 185
rect 674 190 678 201
rect 681 199 685 209
rect 681 197 682 199
rect 684 197 685 199
rect 681 195 685 197
rect 674 189 692 190
rect 654 187 658 189
rect 674 188 688 189
rect 654 185 655 187
rect 657 185 658 187
rect 639 180 649 181
rect 639 178 645 180
rect 647 178 649 180
rect 639 177 649 178
rect 654 180 658 185
rect 663 187 688 188
rect 690 187 692 189
rect 663 185 665 187
rect 667 186 692 187
rect 667 185 678 186
rect 663 184 678 185
rect 654 178 655 180
rect 657 179 679 180
rect 657 178 675 179
rect 654 177 675 178
rect 677 177 679 179
rect 654 176 679 177
rect 684 176 688 178
rect 484 174 485 176
rect 487 174 488 176
rect 585 174 586 176
rect 588 174 589 176
rect 684 174 685 176
rect 687 174 688 176
rect 426 173 432 174
rect 426 171 428 173
rect 430 171 432 173
rect 484 171 488 174
rect 527 173 533 174
rect 527 171 529 173
rect 531 171 533 173
rect 585 171 589 174
rect 626 173 632 174
rect 626 171 628 173
rect 630 171 632 173
rect 684 171 688 174
rect 31 153 33 155
rect 35 153 37 155
rect 31 152 37 153
rect 89 152 93 155
rect 89 150 90 152
rect 92 150 93 152
rect 59 149 84 150
rect 44 148 54 149
rect 44 146 50 148
rect 52 146 54 148
rect 44 145 54 146
rect 59 148 80 149
rect 59 146 60 148
rect 62 147 80 148
rect 82 147 84 149
rect 89 148 93 150
rect 62 146 84 147
rect 44 141 48 145
rect 28 137 48 141
rect 28 134 32 137
rect 26 132 32 134
rect 26 130 27 132
rect 29 130 32 132
rect 26 128 32 130
rect 28 117 32 128
rect 36 132 40 134
rect 59 141 63 146
rect 59 139 60 141
rect 62 139 63 141
rect 59 137 63 139
rect 68 141 83 142
rect 68 139 70 141
rect 72 140 83 141
rect 72 139 97 140
rect 68 138 93 139
rect 79 137 93 138
rect 95 137 97 139
rect 79 136 97 137
rect 36 130 37 132
rect 39 130 40 132
rect 36 125 40 130
rect 79 125 83 136
rect 76 121 83 125
rect 86 129 90 131
rect 86 127 87 129
rect 89 127 90 129
rect 76 120 80 121
rect 76 118 77 120
rect 79 118 80 120
rect 28 116 68 117
rect 76 116 80 118
rect 86 117 90 127
rect 28 114 42 116
rect 44 114 68 116
rect 28 113 68 114
rect 84 113 90 117
rect 41 109 45 113
rect 64 109 88 113
rect 30 108 36 109
rect 30 106 32 108
rect 34 106 36 108
rect 30 101 36 106
rect 41 107 42 109
rect 44 107 45 109
rect 41 105 45 107
rect 52 108 58 109
rect 52 106 54 108
rect 56 106 58 108
rect 30 99 32 101
rect 34 99 36 101
rect 52 101 58 106
rect 118 148 124 155
rect 118 146 120 148
rect 122 146 124 148
rect 118 145 124 146
rect 129 146 133 148
rect 129 144 130 146
rect 132 144 133 146
rect 129 142 133 144
rect 138 146 144 155
rect 172 153 174 155
rect 176 153 178 155
rect 172 152 178 153
rect 230 152 234 155
rect 230 150 231 152
rect 233 150 234 152
rect 272 152 276 155
rect 328 153 330 155
rect 332 153 334 155
rect 328 152 334 153
rect 272 150 273 152
rect 275 150 276 152
rect 200 149 225 150
rect 138 144 140 146
rect 142 144 144 146
rect 138 143 144 144
rect 185 148 195 149
rect 185 146 191 148
rect 193 146 195 148
rect 185 145 195 146
rect 200 148 221 149
rect 200 146 201 148
rect 203 147 221 148
rect 223 147 225 149
rect 230 148 234 150
rect 203 146 225 147
rect 116 138 133 142
rect 116 132 120 138
rect 185 141 189 145
rect 169 137 189 141
rect 169 134 173 137
rect 116 130 117 132
rect 119 130 120 132
rect 116 117 120 130
rect 139 118 140 134
rect 112 110 113 116
rect 116 113 128 117
rect 124 108 128 113
rect 167 132 173 134
rect 167 130 168 132
rect 170 130 173 132
rect 167 128 173 130
rect 169 117 173 128
rect 177 132 181 134
rect 200 141 204 146
rect 200 139 201 141
rect 203 139 204 141
rect 200 137 204 139
rect 209 141 224 142
rect 209 139 211 141
rect 213 140 224 141
rect 213 139 238 140
rect 209 138 234 139
rect 220 137 234 138
rect 236 137 238 139
rect 220 136 238 137
rect 177 130 178 132
rect 180 130 181 132
rect 177 125 181 130
rect 220 125 224 136
rect 217 121 224 125
rect 227 129 231 131
rect 227 127 228 129
rect 230 127 231 129
rect 217 120 221 121
rect 217 118 218 120
rect 220 118 221 120
rect 169 116 209 117
rect 217 116 221 118
rect 227 117 231 127
rect 169 114 183 116
rect 185 114 209 116
rect 169 113 209 114
rect 225 113 231 117
rect 182 109 186 113
rect 205 109 229 113
rect 171 108 177 109
rect 124 107 144 108
rect 124 105 140 107
rect 142 105 144 107
rect 124 104 144 105
rect 171 106 173 108
rect 175 106 177 108
rect 52 99 54 101
rect 56 99 58 101
rect 87 101 93 102
rect 87 99 89 101
rect 91 99 93 101
rect 171 101 177 106
rect 182 107 183 109
rect 185 107 186 109
rect 182 105 186 107
rect 193 108 199 109
rect 193 106 195 108
rect 197 106 199 108
rect 171 99 173 101
rect 175 99 177 101
rect 193 101 199 106
rect 272 148 276 150
rect 281 149 306 150
rect 281 147 283 149
rect 285 148 306 149
rect 285 147 303 148
rect 281 146 303 147
rect 305 146 306 148
rect 282 141 297 142
rect 282 140 293 141
rect 268 139 293 140
rect 295 139 297 141
rect 268 137 270 139
rect 272 138 297 139
rect 302 141 306 146
rect 311 148 321 149
rect 311 146 313 148
rect 315 146 321 148
rect 311 145 321 146
rect 302 139 303 141
rect 305 139 306 141
rect 272 137 286 138
rect 302 137 306 139
rect 268 136 286 137
rect 275 129 279 131
rect 275 127 276 129
rect 278 127 279 129
rect 275 117 279 127
rect 282 125 286 136
rect 317 141 321 145
rect 317 137 337 141
rect 333 134 337 137
rect 325 132 329 134
rect 325 130 326 132
rect 328 130 329 132
rect 325 125 329 130
rect 333 132 339 134
rect 333 130 336 132
rect 338 130 339 132
rect 333 128 339 130
rect 282 121 289 125
rect 285 120 289 121
rect 285 118 286 120
rect 288 118 289 120
rect 275 113 281 117
rect 285 116 289 118
rect 333 117 337 128
rect 297 116 337 117
rect 297 114 321 116
rect 323 114 337 116
rect 297 113 337 114
rect 277 109 301 113
rect 320 109 324 113
rect 372 148 378 155
rect 372 146 374 148
rect 376 146 378 148
rect 372 145 378 146
rect 383 146 387 148
rect 383 144 384 146
rect 386 144 387 146
rect 383 142 387 144
rect 392 146 398 155
rect 426 153 428 155
rect 430 153 432 155
rect 426 152 432 153
rect 484 152 488 155
rect 527 153 529 155
rect 531 153 533 155
rect 527 152 533 153
rect 585 152 589 155
rect 626 153 628 155
rect 630 153 632 155
rect 626 152 632 153
rect 684 152 688 155
rect 484 150 485 152
rect 487 150 488 152
rect 585 150 586 152
rect 588 150 589 152
rect 684 150 685 152
rect 687 150 688 152
rect 454 149 479 150
rect 392 144 394 146
rect 396 144 398 146
rect 392 143 398 144
rect 439 148 449 149
rect 439 146 445 148
rect 447 146 449 148
rect 439 145 449 146
rect 454 148 475 149
rect 454 146 455 148
rect 457 147 475 148
rect 477 147 479 149
rect 484 148 488 150
rect 555 149 580 150
rect 457 146 479 147
rect 370 138 387 142
rect 370 132 374 138
rect 370 130 371 132
rect 373 130 374 132
rect 370 117 374 130
rect 393 118 394 134
rect 366 110 367 116
rect 370 113 382 117
rect 307 108 313 109
rect 307 106 309 108
rect 311 106 313 108
rect 193 99 195 101
rect 197 99 199 101
rect 228 101 234 102
rect 228 99 230 101
rect 232 99 234 101
rect 272 101 278 102
rect 272 99 274 101
rect 276 99 278 101
rect 307 101 313 106
rect 320 107 321 109
rect 323 107 324 109
rect 320 105 324 107
rect 329 108 335 109
rect 329 106 331 108
rect 333 106 335 108
rect 307 99 309 101
rect 311 99 313 101
rect 329 101 335 106
rect 378 108 382 113
rect 439 141 443 145
rect 423 137 443 141
rect 423 134 427 137
rect 421 132 427 134
rect 421 130 422 132
rect 424 130 427 132
rect 421 128 427 130
rect 423 117 427 128
rect 431 132 435 134
rect 454 141 458 146
rect 454 139 455 141
rect 457 139 458 141
rect 454 137 458 139
rect 463 141 478 142
rect 463 139 465 141
rect 467 140 478 141
rect 467 139 492 140
rect 463 138 488 139
rect 474 137 488 138
rect 490 137 492 139
rect 474 136 492 137
rect 431 130 432 132
rect 434 130 435 132
rect 431 125 435 130
rect 474 125 478 136
rect 471 121 478 125
rect 481 129 485 131
rect 481 127 482 129
rect 484 127 485 129
rect 471 120 475 121
rect 471 118 472 120
rect 474 118 475 120
rect 423 116 463 117
rect 471 116 475 118
rect 481 117 485 127
rect 423 114 437 116
rect 439 114 463 116
rect 423 113 463 114
rect 479 113 485 117
rect 436 109 440 113
rect 459 109 483 113
rect 540 148 550 149
rect 540 146 546 148
rect 548 146 550 148
rect 540 145 550 146
rect 555 148 576 149
rect 555 146 556 148
rect 558 147 576 148
rect 578 147 580 149
rect 585 148 589 150
rect 654 149 679 150
rect 558 146 580 147
rect 540 141 544 145
rect 524 137 544 141
rect 524 134 528 137
rect 522 132 528 134
rect 522 130 523 132
rect 525 130 528 132
rect 522 128 528 130
rect 524 117 528 128
rect 532 132 536 134
rect 555 141 559 146
rect 555 139 556 141
rect 558 139 559 141
rect 555 137 559 139
rect 564 141 579 142
rect 564 139 566 141
rect 568 140 579 141
rect 568 139 593 140
rect 564 138 589 139
rect 575 137 589 138
rect 591 137 593 139
rect 575 136 593 137
rect 532 130 533 132
rect 535 130 536 132
rect 532 125 536 130
rect 575 125 579 136
rect 572 121 579 125
rect 582 129 586 131
rect 582 127 583 129
rect 585 127 586 129
rect 572 120 576 121
rect 572 118 573 120
rect 575 118 576 120
rect 524 116 564 117
rect 572 116 576 118
rect 582 117 586 127
rect 524 114 538 116
rect 540 114 564 116
rect 524 113 564 114
rect 580 113 586 117
rect 537 109 541 113
rect 560 109 584 113
rect 639 148 649 149
rect 639 146 645 148
rect 647 146 649 148
rect 639 145 649 146
rect 654 148 675 149
rect 654 146 655 148
rect 657 147 675 148
rect 677 147 679 149
rect 684 148 688 150
rect 657 146 679 147
rect 639 141 643 145
rect 623 137 643 141
rect 623 134 627 137
rect 621 132 627 134
rect 621 130 622 132
rect 624 130 627 132
rect 621 128 627 130
rect 623 117 627 128
rect 631 132 635 134
rect 654 141 658 146
rect 654 139 655 141
rect 657 139 658 141
rect 654 137 658 139
rect 663 141 678 142
rect 663 139 665 141
rect 667 140 678 141
rect 667 139 692 140
rect 663 138 688 139
rect 674 137 688 138
rect 690 137 692 139
rect 674 136 692 137
rect 631 130 632 132
rect 634 130 635 132
rect 631 125 635 130
rect 674 125 678 136
rect 671 121 678 125
rect 681 129 685 131
rect 681 127 682 129
rect 684 127 685 129
rect 671 120 675 121
rect 671 118 672 120
rect 674 118 675 120
rect 623 116 663 117
rect 671 116 675 118
rect 681 117 685 127
rect 623 114 637 116
rect 639 114 663 116
rect 623 113 663 114
rect 679 113 685 117
rect 636 109 640 113
rect 659 109 683 113
rect 425 108 431 109
rect 378 107 398 108
rect 378 105 394 107
rect 396 105 398 107
rect 378 104 398 105
rect 425 106 427 108
rect 429 106 431 108
rect 329 99 331 101
rect 333 99 335 101
rect 425 101 431 106
rect 436 107 437 109
rect 439 107 440 109
rect 436 105 440 107
rect 447 108 453 109
rect 447 106 449 108
rect 451 106 453 108
rect 425 99 427 101
rect 429 99 431 101
rect 447 101 453 106
rect 526 108 532 109
rect 526 106 528 108
rect 530 106 532 108
rect 447 99 449 101
rect 451 99 453 101
rect 482 101 488 102
rect 482 99 484 101
rect 486 99 488 101
rect 526 101 532 106
rect 537 107 538 109
rect 540 107 541 109
rect 537 105 541 107
rect 548 108 554 109
rect 548 106 550 108
rect 552 106 554 108
rect 526 99 528 101
rect 530 99 532 101
rect 548 101 554 106
rect 625 108 631 109
rect 625 106 627 108
rect 629 106 631 108
rect 548 99 550 101
rect 552 99 554 101
rect 583 101 589 102
rect 583 99 585 101
rect 587 99 589 101
rect 625 101 631 106
rect 636 107 637 109
rect 639 107 640 109
rect 636 105 640 107
rect 647 108 653 109
rect 647 106 649 108
rect 651 106 653 108
rect 625 99 627 101
rect 629 99 631 101
rect 647 101 653 106
rect 647 99 649 101
rect 651 99 653 101
rect 682 101 688 102
rect 682 99 684 101
rect 686 99 688 101
rect 69 81 71 83
rect 73 81 75 83
rect 34 77 54 78
rect 34 75 50 77
rect 52 75 54 77
rect 34 74 54 75
rect 69 76 75 81
rect 91 81 93 83
rect 95 81 97 83
rect 69 74 71 76
rect 73 74 75 76
rect 22 66 23 72
rect 34 69 38 74
rect 69 73 75 74
rect 80 75 84 77
rect 80 73 81 75
rect 83 73 84 75
rect 91 76 97 81
rect 126 81 128 83
rect 130 81 132 83
rect 126 80 132 81
rect 170 81 172 83
rect 174 81 176 83
rect 91 74 93 76
rect 95 74 97 76
rect 91 73 97 74
rect 170 76 176 81
rect 192 81 194 83
rect 196 81 198 83
rect 170 74 172 76
rect 174 74 176 76
rect 170 73 176 74
rect 181 75 185 77
rect 181 73 182 75
rect 184 73 185 75
rect 192 76 198 81
rect 227 81 229 83
rect 231 81 233 83
rect 227 80 233 81
rect 271 81 273 83
rect 275 81 277 83
rect 192 74 194 76
rect 196 74 198 76
rect 192 73 198 74
rect 271 76 277 81
rect 293 81 295 83
rect 297 81 299 83
rect 271 74 273 76
rect 275 74 277 76
rect 271 73 277 74
rect 282 75 286 77
rect 282 73 283 75
rect 285 73 286 75
rect 293 76 299 81
rect 328 81 330 83
rect 332 81 334 83
rect 328 80 334 81
rect 424 81 426 83
rect 428 81 430 83
rect 293 74 295 76
rect 297 74 299 76
rect 293 73 299 74
rect 26 65 38 69
rect 80 69 84 73
rect 103 69 127 73
rect 26 52 30 65
rect 26 50 27 52
rect 29 50 30 52
rect 26 44 30 50
rect 49 48 50 64
rect 67 68 107 69
rect 67 66 81 68
rect 83 66 107 68
rect 67 65 107 66
rect 26 40 43 44
rect 39 38 43 40
rect 28 36 34 37
rect 28 34 30 36
rect 32 34 34 36
rect 39 36 40 38
rect 42 36 43 38
rect 39 34 43 36
rect 48 38 54 39
rect 48 36 50 38
rect 52 36 54 38
rect 28 27 34 34
rect 48 27 54 36
rect 67 54 71 65
rect 115 64 119 66
rect 123 65 129 69
rect 115 62 116 64
rect 118 62 119 64
rect 115 61 119 62
rect 115 57 122 61
rect 65 52 71 54
rect 65 50 66 52
rect 68 50 71 52
rect 65 48 71 50
rect 75 52 79 57
rect 75 50 76 52
rect 78 50 79 52
rect 75 48 79 50
rect 67 45 71 48
rect 67 41 87 45
rect 83 37 87 41
rect 118 46 122 57
rect 125 55 129 65
rect 125 53 126 55
rect 128 53 129 55
rect 125 51 129 53
rect 118 45 136 46
rect 98 43 102 45
rect 118 44 132 45
rect 98 41 99 43
rect 101 41 102 43
rect 83 36 93 37
rect 83 34 89 36
rect 91 34 93 36
rect 83 33 93 34
rect 98 36 102 41
rect 107 43 132 44
rect 134 43 136 45
rect 107 41 109 43
rect 111 42 136 43
rect 111 41 122 42
rect 107 40 122 41
rect 98 34 99 36
rect 101 35 123 36
rect 101 34 119 35
rect 98 33 119 34
rect 121 33 123 35
rect 98 32 123 33
rect 128 32 132 34
rect 181 69 185 73
rect 204 69 228 73
rect 168 68 208 69
rect 168 66 182 68
rect 184 66 208 68
rect 168 65 208 66
rect 168 54 172 65
rect 216 64 220 66
rect 224 65 230 69
rect 216 62 217 64
rect 219 62 220 64
rect 216 61 220 62
rect 216 57 223 61
rect 166 52 172 54
rect 166 50 167 52
rect 169 50 172 52
rect 166 48 172 50
rect 176 52 180 57
rect 176 50 177 52
rect 179 50 180 52
rect 176 48 180 50
rect 168 45 172 48
rect 168 41 188 45
rect 184 37 188 41
rect 219 46 223 57
rect 226 55 230 65
rect 226 53 227 55
rect 229 53 230 55
rect 226 51 230 53
rect 219 45 237 46
rect 199 43 203 45
rect 219 44 233 45
rect 199 41 200 43
rect 202 41 203 43
rect 184 36 194 37
rect 184 34 190 36
rect 192 34 194 36
rect 184 33 194 34
rect 199 36 203 41
rect 208 43 233 44
rect 235 43 237 45
rect 208 41 210 43
rect 212 42 237 43
rect 212 41 223 42
rect 208 40 223 41
rect 199 34 200 36
rect 202 35 224 36
rect 202 34 220 35
rect 199 33 220 34
rect 222 33 224 35
rect 199 32 224 33
rect 229 32 233 34
rect 282 69 286 73
rect 305 69 329 73
rect 269 68 309 69
rect 269 66 283 68
rect 285 66 309 68
rect 269 65 309 66
rect 269 54 273 65
rect 317 64 321 66
rect 325 65 331 69
rect 317 62 318 64
rect 320 62 321 64
rect 317 61 321 62
rect 317 57 324 61
rect 267 52 273 54
rect 267 50 268 52
rect 270 50 273 52
rect 267 48 273 50
rect 277 52 281 57
rect 277 50 278 52
rect 280 50 281 52
rect 277 48 281 50
rect 269 45 273 48
rect 269 41 289 45
rect 285 37 289 41
rect 320 46 324 57
rect 327 55 331 65
rect 327 53 328 55
rect 330 53 331 55
rect 327 51 331 53
rect 320 45 338 46
rect 300 43 304 45
rect 320 44 334 45
rect 300 41 301 43
rect 303 41 304 43
rect 285 36 295 37
rect 285 34 291 36
rect 293 34 295 36
rect 285 33 295 34
rect 300 36 304 41
rect 309 43 334 44
rect 336 43 338 45
rect 309 41 311 43
rect 313 42 338 43
rect 313 41 324 42
rect 309 40 324 41
rect 300 34 301 36
rect 303 35 325 36
rect 303 34 321 35
rect 300 33 321 34
rect 323 33 325 35
rect 300 32 325 33
rect 330 32 334 34
rect 377 77 397 78
rect 377 75 393 77
rect 395 75 397 77
rect 377 74 397 75
rect 424 76 430 81
rect 446 81 448 83
rect 450 81 452 83
rect 424 74 426 76
rect 428 74 430 76
rect 365 66 366 72
rect 377 69 381 74
rect 424 73 430 74
rect 435 75 439 77
rect 435 73 436 75
rect 438 73 439 75
rect 446 76 452 81
rect 481 81 483 83
rect 485 81 487 83
rect 481 80 487 81
rect 525 81 527 83
rect 529 81 531 83
rect 446 74 448 76
rect 450 74 452 76
rect 446 73 452 74
rect 525 76 531 81
rect 547 81 549 83
rect 551 81 553 83
rect 525 74 527 76
rect 529 74 531 76
rect 525 73 531 74
rect 536 75 540 77
rect 536 73 537 75
rect 539 73 540 75
rect 547 76 553 81
rect 582 81 584 83
rect 586 81 588 83
rect 582 80 588 81
rect 624 81 626 83
rect 628 81 630 83
rect 547 74 549 76
rect 551 74 553 76
rect 547 73 553 74
rect 624 76 630 81
rect 646 81 648 83
rect 650 81 652 83
rect 624 74 626 76
rect 628 74 630 76
rect 624 73 630 74
rect 635 75 639 77
rect 635 73 636 75
rect 638 73 639 75
rect 646 76 652 81
rect 681 81 683 83
rect 685 81 687 83
rect 681 80 687 81
rect 646 74 648 76
rect 650 74 652 76
rect 646 73 652 74
rect 369 65 381 69
rect 435 69 439 73
rect 458 69 482 73
rect 369 52 373 65
rect 369 50 370 52
rect 372 50 373 52
rect 369 44 373 50
rect 392 48 393 64
rect 422 68 462 69
rect 422 66 436 68
rect 438 66 462 68
rect 422 65 462 66
rect 369 40 386 44
rect 382 38 386 40
rect 371 36 377 37
rect 371 34 373 36
rect 375 34 377 36
rect 382 36 383 38
rect 385 36 386 38
rect 382 34 386 36
rect 391 38 397 39
rect 391 36 393 38
rect 395 36 397 38
rect 128 30 129 32
rect 131 30 132 32
rect 229 30 230 32
rect 232 30 233 32
rect 330 30 331 32
rect 333 30 334 32
rect 70 29 76 30
rect 70 27 72 29
rect 74 27 76 29
rect 128 27 132 30
rect 171 29 177 30
rect 171 27 173 29
rect 175 27 177 29
rect 229 27 233 30
rect 272 29 278 30
rect 272 27 274 29
rect 276 27 278 29
rect 330 27 334 30
rect 371 27 377 34
rect 391 27 397 36
rect 422 54 426 65
rect 470 64 474 66
rect 478 65 484 69
rect 470 62 471 64
rect 473 62 474 64
rect 470 61 474 62
rect 470 57 477 61
rect 420 52 426 54
rect 420 50 421 52
rect 423 50 426 52
rect 420 48 426 50
rect 430 52 434 57
rect 430 50 431 52
rect 433 50 434 52
rect 430 48 434 50
rect 422 45 426 48
rect 422 41 442 45
rect 438 37 442 41
rect 473 46 477 57
rect 480 55 484 65
rect 480 53 481 55
rect 483 53 484 55
rect 480 51 484 53
rect 473 45 491 46
rect 453 43 457 45
rect 473 44 487 45
rect 453 41 454 43
rect 456 41 457 43
rect 438 36 448 37
rect 438 34 444 36
rect 446 34 448 36
rect 438 33 448 34
rect 453 36 457 41
rect 462 43 487 44
rect 489 43 491 45
rect 462 41 464 43
rect 466 42 491 43
rect 466 41 477 42
rect 462 40 477 41
rect 453 34 454 36
rect 456 35 478 36
rect 456 34 474 35
rect 453 33 474 34
rect 476 33 478 35
rect 453 32 478 33
rect 483 32 487 34
rect 536 69 540 73
rect 559 69 583 73
rect 523 68 563 69
rect 523 66 537 68
rect 539 66 563 68
rect 523 65 563 66
rect 523 54 527 65
rect 571 64 575 66
rect 579 65 585 69
rect 571 62 572 64
rect 574 62 575 64
rect 571 61 575 62
rect 571 57 578 61
rect 521 52 527 54
rect 521 50 522 52
rect 524 50 527 52
rect 521 48 527 50
rect 531 52 535 57
rect 531 50 532 52
rect 534 50 535 52
rect 531 48 535 50
rect 523 45 527 48
rect 523 41 543 45
rect 539 37 543 41
rect 574 46 578 57
rect 581 55 585 65
rect 581 53 582 55
rect 584 53 585 55
rect 581 51 585 53
rect 574 45 592 46
rect 554 43 558 45
rect 574 44 588 45
rect 554 41 555 43
rect 557 41 558 43
rect 539 36 549 37
rect 539 34 545 36
rect 547 34 549 36
rect 539 33 549 34
rect 554 36 558 41
rect 563 43 588 44
rect 590 43 592 45
rect 563 41 565 43
rect 567 42 592 43
rect 567 41 578 42
rect 563 40 578 41
rect 554 34 555 36
rect 557 35 579 36
rect 557 34 575 35
rect 554 33 575 34
rect 577 33 579 35
rect 554 32 579 33
rect 584 32 588 34
rect 635 69 639 73
rect 658 69 682 73
rect 622 68 662 69
rect 622 66 636 68
rect 638 66 662 68
rect 622 65 662 66
rect 622 54 626 65
rect 670 64 674 66
rect 678 65 684 69
rect 670 62 671 64
rect 673 62 674 64
rect 670 61 674 62
rect 670 57 677 61
rect 620 52 626 54
rect 620 50 621 52
rect 623 50 626 52
rect 620 48 626 50
rect 630 52 634 57
rect 630 50 631 52
rect 633 50 634 52
rect 630 48 634 50
rect 622 45 626 48
rect 622 41 642 45
rect 638 37 642 41
rect 673 46 677 57
rect 680 55 684 65
rect 680 53 681 55
rect 683 53 684 55
rect 680 51 684 53
rect 673 45 691 46
rect 653 43 657 45
rect 673 44 687 45
rect 653 41 654 43
rect 656 41 657 43
rect 638 36 648 37
rect 638 34 644 36
rect 646 34 648 36
rect 638 33 648 34
rect 653 36 657 41
rect 662 43 687 44
rect 689 43 691 45
rect 662 41 664 43
rect 666 42 691 43
rect 666 41 677 42
rect 662 40 677 41
rect 653 34 654 36
rect 656 35 678 36
rect 656 34 674 35
rect 653 33 674 34
rect 676 33 678 35
rect 653 32 678 33
rect 683 32 687 34
rect 483 30 484 32
rect 486 30 487 32
rect 584 30 585 32
rect 587 30 588 32
rect 683 30 684 32
rect 686 30 687 32
rect 425 29 431 30
rect 425 27 427 29
rect 429 27 431 29
rect 483 27 487 30
rect 526 29 532 30
rect 526 27 528 29
rect 530 27 532 29
rect 584 27 588 30
rect 625 29 631 30
rect 625 27 627 29
rect 629 27 631 29
rect 683 27 687 30
<< via1 >>
rect 50 362 52 364
rect 28 346 30 348
rect 26 329 28 331
rect 59 346 61 348
rect 66 329 68 331
rect 90 321 92 323
rect 115 346 117 348
rect 132 329 134 331
rect 117 322 119 324
rect 179 322 181 324
rect 261 346 263 348
rect 244 329 246 331
rect 197 322 199 324
rect 259 322 261 324
rect 326 362 328 364
rect 317 346 319 348
rect 286 321 288 323
rect 310 329 312 331
rect 348 346 350 348
rect 350 329 352 331
rect 431 346 433 348
rect 414 329 416 331
rect 367 322 369 324
rect 429 322 431 324
rect 496 362 498 364
rect 487 346 489 348
rect 566 362 568 364
rect 456 321 458 323
rect 480 329 482 331
rect 518 346 520 348
rect 544 346 546 348
rect 520 329 522 331
rect 542 329 544 331
rect 575 346 577 348
rect 582 329 584 331
rect 606 321 608 323
rect 631 346 633 348
rect 648 329 650 331
rect 633 322 635 324
rect 26 283 28 285
rect 28 266 30 268
rect 51 274 53 276
rect 66 283 68 285
rect 90 291 92 293
rect 59 266 61 268
rect 123 274 125 276
rect 115 266 117 268
rect 179 255 181 257
rect 253 274 255 276
rect 261 266 263 268
rect 275 258 277 260
rect 197 255 199 257
rect 286 291 288 293
rect 310 283 312 285
rect 317 266 319 268
rect 350 283 352 285
rect 348 266 350 268
rect 326 253 328 255
rect 367 262 369 264
rect 447 282 449 284
rect 423 274 425 276
rect 431 266 433 268
rect 456 291 458 293
rect 480 283 482 285
rect 520 283 522 285
rect 495 274 497 276
rect 487 266 489 268
rect 542 283 544 285
rect 518 266 520 268
rect 544 266 546 268
rect 582 283 584 285
rect 606 291 608 293
rect 575 266 577 268
rect 617 258 619 260
rect 639 274 641 276
rect 631 266 633 268
rect 687 250 689 252
rect 140 218 142 220
rect 40 193 42 195
rect 20 178 22 180
rect 109 202 111 204
rect 92 185 94 187
rect 197 202 199 204
rect 194 194 196 196
rect 162 178 164 180
rect 240 178 242 180
rect 278 202 280 204
rect 295 185 297 187
rect 342 178 344 180
rect 363 194 365 196
rect 386 193 388 195
rect 431 202 433 204
rect 449 194 451 196
rect 492 177 494 179
rect 532 202 534 204
rect 516 185 518 187
rect 597 193 599 195
rect 549 185 551 187
rect 631 202 633 204
rect 639 194 641 196
rect 615 185 617 187
rect 695 178 697 180
rect 38 146 40 148
rect 100 146 102 148
rect 53 138 55 140
rect 70 122 72 124
rect 110 139 112 141
rect 194 139 196 141
rect 132 131 134 133
rect 242 138 244 140
rect 214 130 216 132
rect 325 146 327 148
rect 310 138 312 140
rect 327 122 329 124
rect 363 122 365 124
rect 386 131 388 133
rect 271 106 273 108
rect 449 130 451 132
rect 465 122 467 124
rect 516 139 518 141
rect 549 139 551 141
rect 597 131 599 133
rect 566 123 568 125
rect 615 139 617 141
rect 648 139 650 141
rect 665 122 667 124
rect 42 49 44 51
rect 75 58 77 60
rect 93 50 95 52
rect 176 58 178 60
rect 160 41 162 43
rect 241 49 243 51
rect 193 41 195 43
rect 277 58 279 60
rect 261 41 263 43
rect 294 46 296 48
rect 362 46 364 48
rect 385 49 387 51
rect 430 58 432 60
rect 448 50 450 52
rect 531 58 533 60
rect 515 41 517 43
rect 596 49 598 51
rect 548 41 550 43
rect 630 58 632 60
rect 638 50 640 52
rect 614 41 616 43
<< via2 >>
rect 348 370 350 372
rect 544 370 546 372
rect 115 362 117 364
rect 261 362 263 364
rect 431 362 433 364
rect 631 362 633 364
rect 59 354 61 356
rect 487 354 489 356
rect 59 346 61 348
rect 115 346 117 348
rect 261 346 263 348
rect 348 346 350 348
rect 431 346 433 348
rect 487 346 489 348
rect 544 346 546 348
rect 631 346 633 348
rect 26 338 28 340
rect 350 338 352 340
rect 480 337 482 339
rect 582 337 584 339
rect 26 329 28 331
rect 66 329 68 331
rect 132 329 134 331
rect 244 329 246 331
rect 310 329 312 331
rect 350 329 352 331
rect 414 329 416 331
rect 480 329 482 331
rect 520 329 522 331
rect 542 329 544 331
rect 582 329 584 331
rect 648 329 650 331
rect 94 321 96 323
rect 117 322 119 324
rect 184 322 186 324
rect 197 322 199 324
rect 259 322 261 324
rect 282 321 284 323
rect 367 322 369 324
rect 429 322 431 324
rect 452 321 454 323
rect 610 321 612 323
rect 633 322 635 324
rect 132 291 134 293
rect 244 291 246 293
rect 414 291 416 293
rect 648 291 650 293
rect 26 283 28 285
rect 66 283 68 285
rect 310 283 312 285
rect 350 283 352 285
rect 406 282 408 284
rect 480 283 482 285
rect 520 283 522 285
rect 542 283 544 285
rect 582 283 584 285
rect 47 274 49 276
rect 117 274 119 276
rect 196 274 198 276
rect 245 274 247 276
rect 259 274 261 276
rect 429 274 431 276
rect 506 274 508 276
rect 633 274 635 276
rect 55 266 57 268
rect 94 266 96 268
rect 156 266 158 268
rect 206 266 208 268
rect 282 266 284 268
rect 348 266 350 268
rect 452 266 454 268
rect 487 266 489 268
rect 544 266 546 268
rect 610 266 612 268
rect 357 262 359 264
rect 101 258 103 260
rect 206 258 208 260
rect 175 255 177 257
rect 601 258 603 260
rect 197 255 199 257
rect 326 253 328 255
rect 348 253 350 255
rect 544 253 546 255
rect 687 250 689 252
rect 55 245 57 247
rect 487 245 489 247
rect 278 218 280 220
rect 326 218 328 220
rect 631 218 633 220
rect 245 210 247 212
rect 431 210 433 212
rect 506 210 508 212
rect 639 210 641 212
rect 148 202 150 204
rect 197 202 199 204
rect 278 202 280 204
rect 306 202 308 204
rect 406 202 408 204
rect 431 202 433 204
rect 532 202 534 204
rect 631 202 633 204
rect 40 193 42 195
rect 101 193 103 195
rect 109 193 111 195
rect 639 194 641 196
rect 100 185 102 187
rect 148 186 150 188
rect 252 186 254 188
rect 295 185 297 187
rect 20 178 22 180
rect 132 178 134 180
rect 194 178 196 180
rect 252 177 254 179
rect 306 177 308 179
rect 342 178 344 180
rect 492 177 494 179
rect 648 178 650 180
rect 367 169 369 171
rect 532 169 534 171
rect 38 146 40 148
rect 100 146 102 148
rect 295 146 297 148
rect 194 139 196 141
rect 648 139 650 141
rect 132 131 134 133
rect 357 130 359 132
rect 156 122 158 124
rect 492 122 494 124
rect 601 123 603 125
rect 687 122 689 124
rect 271 106 273 108
rect 271 98 273 100
rect 638 98 640 100
rect 342 80 344 82
rect 430 80 432 82
rect 175 66 177 68
rect 277 66 279 68
rect 20 58 22 60
rect 109 58 111 60
rect 277 58 279 60
rect 430 58 432 60
rect 531 58 533 60
rect 630 58 632 60
rect 638 50 640 52
rect 184 33 186 35
rect 531 33 533 35
rect 48 25 50 27
rect 630 25 632 27
<< labels >>
rlabel alu1 100 274 100 274 1 p3
rlabel alu1 101 263 101 263 1 p3
rlabel alu1 173 251 173 251 1 p2
rlabel alu1 181 275 181 275 1 p2
rlabel alu1 173 363 173 363 1 p1
rlabel alu1 181 339 181 339 1 p1
rlabel alu1 137 375 137 375 4 vdd
rlabel alu1 137 311 137 311 4 vss
rlabel alu1 137 303 137 303 2 vss
rlabel alu1 68 267 68 267 1 b2
rlabel alu1 60 259 60 259 1 b2
rlabel alu1 76 339 76 339 1 a3
rlabel alu1 68 335 68 335 1 a3
rlabel alu1 68 347 68 347 1 b3
rlabel alu1 60 355 60 355 1 b3
rlabel alu1 76 303 76 303 2 vss
rlabel alu1 76 375 76 375 4 vdd
rlabel alu1 76 311 76 311 4 vss
rlabel alu1 52 271 52 271 1 p0
rlabel alu1 44 291 44 291 1 p0
rlabel alu1 20 355 20 355 1 b3
rlabel alu1 28 347 28 347 1 b3
rlabel alu1 36 339 36 339 1 a2
rlabel alu1 28 335 28 335 1 a2
rlabel alu1 20 259 20 259 1 b2
rlabel alu1 28 267 28 267 1 b2
rlabel alu1 36 275 36 275 1 a2
rlabel alu1 28 279 28 279 1 a2
rlabel alu1 36 303 36 303 2 vss
rlabel alu1 36 375 36 375 4 vdd
rlabel alu1 36 311 36 311 4 vss
rlabel alu1 67 279 67 279 1 a3
rlabel alu1 310 279 310 279 1 a3
rlabel alu1 310 335 310 335 1 a3
rlabel alu1 310 347 310 347 1 b1
rlabel alu1 318 355 318 355 1 b1
rlabel alu1 358 355 358 355 1 b1
rlabel via1 350 347 350 347 1 b1
rlabel alu1 318 259 318 259 1 b0
rlabel alu1 310 267 310 267 1 b0
rlabel via1 350 267 350 267 1 b0
rlabel alu1 358 259 358 259 1 b0
rlabel alu1 205 363 205 363 1 q1
rlabel alu1 197 339 197 339 1 q1
rlabel alu1 205 251 205 251 1 q2
rlabel alu1 197 275 197 275 1 q2
rlabel alu1 277 263 277 263 1 q3
rlabel alu1 278 274 278 274 1 q3
rlabel alu1 326 271 326 271 1 q0
rlabel alu1 334 291 334 291 1 q0
rlabel alu1 241 375 241 375 6 vdd
rlabel alu1 241 311 241 311 6 vss
rlabel alu1 241 303 241 303 8 vss
rlabel alu1 302 339 302 339 1 a3
rlabel alu1 302 303 302 303 8 vss
rlabel alu1 302 375 302 375 6 vdd
rlabel alu1 302 311 302 311 6 vss
rlabel alu1 342 339 342 339 1 a2
rlabel alu1 350 335 350 335 1 a2
rlabel alu1 342 275 342 275 1 a2
rlabel alu1 350 279 350 279 1 a2
rlabel alu1 342 303 342 303 8 vss
rlabel alu1 342 375 342 375 6 vdd
rlabel alu1 342 311 342 311 6 vss
rlabel alu1 480 279 480 279 1 a1
rlabel alu1 472 339 472 339 1 a1
rlabel alu1 480 335 480 335 1 a1
rlabel alu1 512 339 512 339 1 a0
rlabel alu1 520 335 520 335 1 a0
rlabel alu1 520 279 520 279 1 a0
rlabel alu1 512 275 512 275 1 a0
rlabel alu1 375 363 375 363 1 r1
rlabel alu1 367 339 367 339 1 r1
rlabel alu1 367 275 367 275 1 r2
rlabel alu1 375 251 375 251 1 r2
rlabel alu1 448 274 448 274 1 r3
rlabel alu1 447 263 447 263 1 r3
rlabel alu1 504 291 504 291 1 r0
rlabel alu1 496 271 496 271 1 r0
rlabel alu1 411 375 411 375 6 vdd
rlabel alu1 411 311 411 311 6 vss
rlabel alu1 411 303 411 303 8 vss
rlabel alu1 480 267 480 267 1 b2
rlabel alu1 488 259 488 259 1 b2
rlabel alu1 480 347 480 347 1 b3
rlabel alu1 488 355 488 355 1 b3
rlabel alu1 472 303 472 303 8 vss
rlabel alu1 472 375 472 375 6 vdd
rlabel alu1 472 311 472 311 6 vss
rlabel alu1 528 355 528 355 1 b3
rlabel alu1 520 347 520 347 1 b3
rlabel alu1 528 259 528 259 1 b2
rlabel alu1 520 267 520 267 1 b2
rlabel alu1 512 303 512 303 8 vss
rlabel alu1 512 375 512 375 6 vdd
rlabel alu1 512 311 512 311 6 vss
rlabel alu1 583 279 583 279 1 a1
rlabel alu1 592 339 592 339 1 a1
rlabel alu1 584 335 584 335 1 a1
rlabel alu1 584 347 584 347 1 b1
rlabel alu1 576 355 576 355 1 b1
rlabel alu1 536 355 536 355 1 b1
rlabel via1 544 347 544 347 1 b1
rlabel alu1 552 339 552 339 1 a0
rlabel alu1 544 335 544 335 1 a0
rlabel alu1 584 267 584 267 1 b0
rlabel alu1 576 259 576 259 1 b0
rlabel via1 544 267 544 267 1 b0
rlabel alu1 536 259 536 259 1 b0
rlabel alu1 544 279 544 279 1 a0
rlabel alu1 552 275 552 275 1 a0
rlabel alu1 689 363 689 363 1 o1
rlabel alu1 697 339 697 339 1 o1
rlabel alu1 689 251 689 251 1 s2
rlabel alu1 616 274 616 274 1 s3
rlabel alu1 617 263 617 263 1 s3
rlabel alu1 560 291 560 291 1 o0
rlabel alu1 568 271 568 271 1 o0
rlabel alu1 653 375 653 375 4 vdd
rlabel alu1 653 311 653 311 4 vss
rlabel alu1 653 303 653 303 2 vss
rlabel alu1 592 303 592 303 2 vss
rlabel alu1 592 375 592 375 4 vdd
rlabel alu1 592 311 592 311 4 vss
rlabel alu1 552 303 552 303 2 vss
rlabel alu1 552 375 552 375 4 vdd
rlabel alu1 552 311 552 311 4 vss
rlabel alu1 697 275 697 275 1 s2
rlabel alu1 696 54 696 54 1 o4
rlabel alu1 648 59 648 59 1 p0
rlabel alu1 648 47 648 47 1 u0
rlabel alu1 652 87 652 87 4 vdd
rlabel alu1 652 23 652 23 4 vss
rlabel alu1 653 167 653 167 4 vss
rlabel alu1 653 231 653 231 4 vdd
rlabel alu1 649 191 649 191 1 r0
rlabel alu1 641 195 641 195 1 r0
rlabel pmos 633 203 633 203 1 q0
rlabel alu1 641 203 641 203 1 q0
rlabel alu1 649 203 649 203 1 q0
rlabel alu1 657 203 657 203 1 q0
rlabel alu1 665 199 665 199 1 q0
rlabel alu1 653 159 653 159 2 vss
rlabel alu1 653 95 653 95 2 vdd
rlabel alu1 648 123 648 123 1 s2
rlabel alu1 658 123 658 123 1 s2
rlabel alu1 697 198 697 198 1 t5
rlabel alu1 616 132 616 132 1 t4
rlabel alu1 616 198 616 198 1 t3
rlabel alu1 628 179 628 179 1 t3
rlabel alu1 697 132 697 132 1 o2
rlabel alu1 552 123 552 123 1 s3
rlabel alu1 554 159 554 159 2 vss
rlabel alu1 554 95 554 95 2 vdd
rlabel pmos 534 203 534 203 1 r1
rlabel alu1 542 203 542 203 1 r1
rlabel alu1 550 203 550 203 1 r1
rlabel alu1 558 203 558 203 1 r1
rlabel alu1 566 199 566 199 1 r1
rlabel alu1 554 167 554 167 4 vss
rlabel alu1 554 231 554 231 4 vdd
rlabel alu1 553 87 553 87 4 vdd
rlabel alu1 553 23 553 23 4 vss
rlabel alu1 548 59 548 59 1 p1
rlabel alu1 497 124 497 124 1 o3
rlabel alu1 497 198 497 198 1 t6
rlabel alu1 453 159 453 159 2 vss
rlabel alu1 453 95 453 95 2 vdd
rlabel alu1 465 199 465 199 1 q1
rlabel alu1 457 203 457 203 1 q1
rlabel alu1 449 203 449 203 1 q1
rlabel alu1 441 203 441 203 1 q1
rlabel pmos 433 203 433 203 1 q1
rlabel alu1 453 167 453 167 4 vss
rlabel alu1 453 231 453 231 4 vdd
rlabel alu1 452 87 452 87 4 vdd
rlabel alu1 452 23 452 23 4 vss
rlabel alu1 449 59 449 59 1 u1
rlabel alu1 496 56 496 56 1 o5
rlabel alu1 364 126 364 126 1 t2
rlabel alu1 364 198 364 198 1 t1
rlabel alu1 380 95 380 95 8 vdd
rlabel alu1 380 159 380 159 8 vss
rlabel alu1 380 231 380 231 6 vdd
rlabel alu1 380 167 380 167 6 vss
rlabel alu1 379 23 379 23 6 vss
rlabel alu1 379 87 379 87 6 vdd
rlabel alu1 344 189 344 189 1 u1
rlabel alu1 263 124 263 124 1 u0
rlabel alu1 300 231 300 231 4 vdd
rlabel alu1 300 167 300 167 4 vss
rlabel alu1 307 95 307 95 8 vdd
rlabel alu1 307 159 307 159 8 vss
rlabel alu1 343 55 343 55 1 o6
rlabel alu1 295 59 295 59 1 p2
rlabel alu1 299 87 299 87 4 vdd
rlabel alu1 299 23 299 23 4 vss
rlabel alu1 203 123 203 123 1 r2
rlabel alu1 195 123 195 123 1 r2
rlabel alu1 187 123 187 123 1 r2
rlabel pmos 179 123 179 123 1 r2
rlabel alu1 210 199 210 199 1 q2
rlabel alu1 202 203 202 203 1 q2
rlabel alu1 194 203 194 203 1 q2
rlabel alu1 186 203 186 203 1 q2
rlabel pmos 178 203 178 203 1 q2
rlabel alu1 198 167 198 167 4 vss
rlabel alu1 198 231 198 231 4 vdd
rlabel alu1 199 95 199 95 2 vdd
rlabel alu1 199 159 199 159 2 vss
rlabel alu1 195 59 195 59 1 p3
rlabel alu1 198 23 198 23 4 vss
rlabel alu1 198 87 198 87 4 vdd
rlabel alu1 20 199 20 199 1 ca1
rlabel alu1 109 199 109 199 1 r3
rlabel alu1 101 203 101 203 1 r3
rlabel alu1 93 203 93 203 1 r3
rlabel alu1 85 203 85 203 1 r3
rlabel pmos 77 203 77 203 1 r3
rlabel alu1 62 123 62 123 1 q3
rlabel alu1 54 123 54 123 1 q3
rlabel alu1 46 123 46 123 1 q3
rlabel pmos 38 123 38 123 1 q3
rlabel alu1 126 95 126 95 8 vdd
rlabel alu1 126 159 126 159 8 vss
rlabel alu1 118 107 118 107 8 z
rlabel alu1 110 127 110 127 8 z
rlabel alu1 58 95 58 95 2 vdd
rlabel alu1 58 159 58 159 2 vss
rlabel alu0 69 199 69 199 4 con
rlabel alu1 97 167 97 167 4 vss
rlabel alu1 97 231 97 231 4 vdd
rlabel alu1 36 231 36 231 6 vdd
rlabel alu1 36 167 36 167 6 vss
rlabel alu1 141 55 141 55 1 o7
rlabel alu1 95 59 95 59 1 ca1
rlabel alu1 97 23 97 23 4 vss
rlabel alu1 97 87 97 87 4 vdd
rlabel alu1 36 87 36 87 6 vdd
rlabel alu1 36 23 36 23 6 vss
rlabel alu1 615 47 615 47 1 x1
rlabel alu1 363 56 363 56 1 x2
rlabel alu1 262 52 262 52 1 x3
rlabel alu1 20 53 20 53 1 ca3
<< end >>
