magic
tech scmos
timestamp 1509181223
<< ab >>
rect 69 436 109 580
rect 111 436 238 580
rect 246 436 373 580
rect 375 436 415 580
rect 416 436 543 580
rect 545 436 625 580
rect 627 436 754 580
rect 69 364 453 436
rect 67 360 453 364
rect 64 300 453 360
rect 67 292 453 300
rect 466 292 754 436
rect 69 220 109 292
rect 110 220 452 292
rect 465 220 753 292
<< nwell >>
rect 64 540 758 585
rect 64 396 758 476
rect 64 252 758 332
<< pwell >>
rect 64 476 758 540
rect 64 332 758 396
rect 64 215 758 252
<< poly >>
rect 78 574 80 578
rect 88 574 90 578
rect 98 574 100 578
rect 118 574 120 578
rect 128 574 130 578
rect 138 574 140 578
rect 159 574 161 578
rect 169 574 171 578
rect 179 574 181 578
rect 78 551 80 555
rect 74 549 80 551
rect 74 547 76 549
rect 78 547 80 549
rect 74 545 80 547
rect 78 534 80 545
rect 88 543 90 555
rect 118 551 120 555
rect 114 549 120 551
rect 114 547 116 549
rect 118 547 120 549
rect 98 543 100 546
rect 114 545 120 547
rect 84 541 90 543
rect 84 539 86 541
rect 88 539 90 541
rect 84 537 90 539
rect 94 541 100 543
rect 94 539 96 541
rect 98 539 100 541
rect 94 537 100 539
rect 85 534 87 537
rect 98 534 100 537
rect 118 534 120 545
rect 128 543 130 555
rect 197 571 199 576
rect 204 571 206 576
rect 227 574 229 578
rect 255 574 257 578
rect 214 562 216 567
rect 278 571 280 576
rect 285 571 287 576
rect 303 574 305 578
rect 313 574 315 578
rect 323 574 325 578
rect 344 574 346 578
rect 354 574 356 578
rect 364 574 366 578
rect 384 574 386 578
rect 394 574 396 578
rect 404 574 406 578
rect 425 574 427 578
rect 268 562 270 567
rect 214 546 216 549
rect 138 543 140 546
rect 159 543 161 546
rect 169 543 171 546
rect 179 543 181 546
rect 197 543 199 546
rect 204 543 206 546
rect 214 544 223 546
rect 124 541 130 543
rect 124 539 126 541
rect 128 539 130 541
rect 124 537 130 539
rect 134 541 140 543
rect 134 539 136 541
rect 138 539 140 541
rect 134 537 140 539
rect 157 541 163 543
rect 157 539 159 541
rect 161 539 163 541
rect 157 537 163 539
rect 167 541 173 543
rect 167 539 169 541
rect 171 539 173 541
rect 167 537 173 539
rect 177 541 199 543
rect 177 539 179 541
rect 181 539 186 541
rect 188 539 199 541
rect 177 537 199 539
rect 203 541 209 543
rect 203 539 205 541
rect 207 539 209 541
rect 203 537 209 539
rect 125 534 127 537
rect 138 534 140 537
rect 78 516 80 521
rect 85 516 87 521
rect 98 515 100 520
rect 118 516 120 521
rect 125 516 127 521
rect 159 528 161 537
rect 170 534 172 537
rect 177 534 179 537
rect 197 534 199 537
rect 207 534 209 537
rect 217 542 219 544
rect 221 542 223 544
rect 217 540 223 542
rect 138 515 140 520
rect 217 527 219 540
rect 227 536 229 549
rect 223 534 229 536
rect 223 532 225 534
rect 227 532 229 534
rect 223 530 229 532
rect 227 527 229 530
rect 255 536 257 549
rect 268 546 270 549
rect 261 544 270 546
rect 261 542 263 544
rect 265 542 267 544
rect 278 543 280 546
rect 285 543 287 546
rect 303 543 305 546
rect 313 543 315 546
rect 323 543 325 546
rect 344 543 346 546
rect 354 543 356 555
rect 364 551 366 555
rect 364 549 370 551
rect 364 547 366 549
rect 368 547 370 549
rect 364 545 370 547
rect 261 540 267 542
rect 255 534 261 536
rect 255 532 257 534
rect 259 532 261 534
rect 255 530 261 532
rect 255 527 257 530
rect 265 527 267 540
rect 275 541 281 543
rect 275 539 277 541
rect 279 539 281 541
rect 275 537 281 539
rect 285 541 307 543
rect 285 539 296 541
rect 298 539 303 541
rect 305 539 307 541
rect 285 537 307 539
rect 311 541 317 543
rect 311 539 313 541
rect 315 539 317 541
rect 311 537 317 539
rect 321 541 327 543
rect 321 539 323 541
rect 325 539 327 541
rect 321 537 327 539
rect 344 541 350 543
rect 344 539 346 541
rect 348 539 350 541
rect 344 537 350 539
rect 354 541 360 543
rect 354 539 356 541
rect 358 539 360 541
rect 354 537 360 539
rect 275 534 277 537
rect 285 534 287 537
rect 305 534 307 537
rect 312 534 314 537
rect 197 515 199 520
rect 207 515 209 520
rect 159 510 161 514
rect 170 510 172 514
rect 177 510 179 514
rect 217 512 219 517
rect 227 510 229 514
rect 255 510 257 514
rect 265 512 267 517
rect 275 515 277 520
rect 285 515 287 520
rect 323 528 325 537
rect 344 534 346 537
rect 357 534 359 537
rect 364 534 366 545
rect 384 543 386 546
rect 394 543 396 555
rect 404 551 406 555
rect 404 549 410 551
rect 448 571 450 576
rect 455 571 457 576
rect 473 574 475 578
rect 483 574 485 578
rect 493 574 495 578
rect 514 574 516 578
rect 524 574 526 578
rect 534 574 536 578
rect 554 574 556 578
rect 564 574 566 578
rect 574 574 576 578
rect 594 574 596 578
rect 604 574 606 578
rect 614 574 616 578
rect 634 574 636 578
rect 644 574 646 578
rect 654 574 656 578
rect 675 574 677 578
rect 685 574 687 578
rect 695 574 697 578
rect 438 562 440 567
rect 404 547 406 549
rect 408 547 410 549
rect 404 545 410 547
rect 384 541 390 543
rect 384 539 386 541
rect 388 539 390 541
rect 384 537 390 539
rect 394 541 400 543
rect 394 539 396 541
rect 398 539 400 541
rect 394 537 400 539
rect 384 534 386 537
rect 397 534 399 537
rect 404 534 406 545
rect 425 536 427 549
rect 438 546 440 549
rect 431 544 440 546
rect 431 542 433 544
rect 435 542 437 544
rect 448 543 450 546
rect 455 543 457 546
rect 473 543 475 546
rect 483 543 485 546
rect 493 543 495 546
rect 514 543 516 546
rect 524 543 526 555
rect 534 551 536 555
rect 534 549 540 551
rect 534 547 536 549
rect 538 547 540 549
rect 534 545 540 547
rect 431 540 437 542
rect 425 534 431 536
rect 344 515 346 520
rect 357 516 359 521
rect 364 516 366 521
rect 425 532 427 534
rect 429 532 431 534
rect 425 530 431 532
rect 425 527 427 530
rect 435 527 437 540
rect 445 541 451 543
rect 445 539 447 541
rect 449 539 451 541
rect 445 537 451 539
rect 455 541 477 543
rect 455 539 466 541
rect 468 539 473 541
rect 475 539 477 541
rect 455 537 477 539
rect 481 541 487 543
rect 481 539 483 541
rect 485 539 487 541
rect 481 537 487 539
rect 491 541 497 543
rect 491 539 493 541
rect 495 539 497 541
rect 491 537 497 539
rect 514 541 520 543
rect 514 539 516 541
rect 518 539 520 541
rect 514 537 520 539
rect 524 541 530 543
rect 524 539 526 541
rect 528 539 530 541
rect 524 537 530 539
rect 445 534 447 537
rect 455 534 457 537
rect 475 534 477 537
rect 482 534 484 537
rect 384 515 386 520
rect 397 516 399 521
rect 404 516 406 521
rect 305 510 307 514
rect 312 510 314 514
rect 323 510 325 514
rect 425 510 427 514
rect 435 512 437 517
rect 445 515 447 520
rect 455 515 457 520
rect 493 528 495 537
rect 514 534 516 537
rect 527 534 529 537
rect 534 534 536 545
rect 554 543 556 546
rect 564 543 566 555
rect 574 551 576 555
rect 594 551 596 555
rect 574 549 580 551
rect 574 547 576 549
rect 578 547 580 549
rect 574 545 580 547
rect 590 549 596 551
rect 590 547 592 549
rect 594 547 596 549
rect 590 545 596 547
rect 554 541 560 543
rect 554 539 556 541
rect 558 539 560 541
rect 554 537 560 539
rect 564 541 570 543
rect 564 539 566 541
rect 568 539 570 541
rect 564 537 570 539
rect 554 534 556 537
rect 567 534 569 537
rect 574 534 576 545
rect 594 534 596 545
rect 604 543 606 555
rect 634 551 636 555
rect 630 549 636 551
rect 630 547 632 549
rect 634 547 636 549
rect 614 543 616 546
rect 630 545 636 547
rect 600 541 606 543
rect 600 539 602 541
rect 604 539 606 541
rect 600 537 606 539
rect 610 541 616 543
rect 610 539 612 541
rect 614 539 616 541
rect 610 537 616 539
rect 601 534 603 537
rect 614 534 616 537
rect 634 534 636 545
rect 644 543 646 555
rect 713 571 715 576
rect 720 571 722 576
rect 743 574 745 578
rect 730 562 732 567
rect 730 546 732 549
rect 654 543 656 546
rect 675 543 677 546
rect 685 543 687 546
rect 695 543 697 546
rect 713 543 715 546
rect 720 543 722 546
rect 730 544 739 546
rect 640 541 646 543
rect 640 539 642 541
rect 644 539 646 541
rect 640 537 646 539
rect 650 541 656 543
rect 650 539 652 541
rect 654 539 656 541
rect 650 537 656 539
rect 673 541 679 543
rect 673 539 675 541
rect 677 539 679 541
rect 673 537 679 539
rect 683 541 689 543
rect 683 539 685 541
rect 687 539 689 541
rect 683 537 689 539
rect 693 541 715 543
rect 693 539 695 541
rect 697 539 702 541
rect 704 539 715 541
rect 693 537 715 539
rect 719 541 725 543
rect 719 539 721 541
rect 723 539 725 541
rect 719 537 725 539
rect 641 534 643 537
rect 654 534 656 537
rect 514 515 516 520
rect 527 516 529 521
rect 534 516 536 521
rect 554 515 556 520
rect 567 516 569 521
rect 574 516 576 521
rect 594 516 596 521
rect 601 516 603 521
rect 475 510 477 514
rect 482 510 484 514
rect 493 510 495 514
rect 614 515 616 520
rect 634 516 636 521
rect 641 516 643 521
rect 675 528 677 537
rect 686 534 688 537
rect 693 534 695 537
rect 713 534 715 537
rect 723 534 725 537
rect 733 542 735 544
rect 737 542 739 544
rect 733 540 739 542
rect 654 515 656 520
rect 733 527 735 540
rect 743 536 745 549
rect 739 534 745 536
rect 739 532 741 534
rect 743 532 745 534
rect 739 530 745 532
rect 743 527 745 530
rect 713 515 715 520
rect 723 515 725 520
rect 675 510 677 514
rect 686 510 688 514
rect 693 510 695 514
rect 733 512 735 517
rect 743 510 745 514
rect 159 502 161 506
rect 170 502 172 506
rect 177 502 179 506
rect 78 495 80 500
rect 85 495 87 500
rect 98 496 100 501
rect 118 495 120 500
rect 125 495 127 500
rect 138 496 140 501
rect 78 471 80 482
rect 85 479 87 482
rect 98 479 100 482
rect 84 477 90 479
rect 84 475 86 477
rect 88 475 90 477
rect 84 473 90 475
rect 94 477 100 479
rect 94 475 96 477
rect 98 475 100 477
rect 94 473 100 475
rect 74 469 80 471
rect 74 467 76 469
rect 78 467 80 469
rect 74 465 80 467
rect 78 461 80 465
rect 88 461 90 473
rect 98 470 100 473
rect 118 471 120 482
rect 125 479 127 482
rect 138 479 140 482
rect 159 479 161 488
rect 197 496 199 501
rect 207 496 209 501
rect 217 499 219 504
rect 227 502 229 506
rect 255 502 257 506
rect 265 499 267 504
rect 305 502 307 506
rect 312 502 314 506
rect 323 502 325 506
rect 275 496 277 501
rect 285 496 287 501
rect 170 479 172 482
rect 177 479 179 482
rect 197 479 199 482
rect 207 479 209 482
rect 124 477 130 479
rect 124 475 126 477
rect 128 475 130 477
rect 124 473 130 475
rect 134 477 140 479
rect 134 475 136 477
rect 138 475 140 477
rect 134 473 140 475
rect 157 477 163 479
rect 157 475 159 477
rect 161 475 163 477
rect 157 473 163 475
rect 167 477 173 479
rect 167 475 169 477
rect 171 475 173 477
rect 167 473 173 475
rect 177 477 199 479
rect 177 475 179 477
rect 181 475 186 477
rect 188 475 199 477
rect 177 473 199 475
rect 203 477 209 479
rect 203 475 205 477
rect 207 475 209 477
rect 203 473 209 475
rect 217 476 219 489
rect 227 486 229 489
rect 223 484 229 486
rect 223 482 225 484
rect 227 482 229 484
rect 223 480 229 482
rect 217 474 223 476
rect 114 469 120 471
rect 114 467 116 469
rect 118 467 120 469
rect 114 465 120 467
rect 118 461 120 465
rect 128 461 130 473
rect 138 470 140 473
rect 159 470 161 473
rect 169 470 171 473
rect 179 470 181 473
rect 197 470 199 473
rect 204 470 206 473
rect 217 472 219 474
rect 221 472 223 474
rect 214 470 223 472
rect 214 467 216 470
rect 227 467 229 480
rect 255 486 257 489
rect 255 484 261 486
rect 255 482 257 484
rect 259 482 261 484
rect 255 480 261 482
rect 255 467 257 480
rect 265 476 267 489
rect 425 502 427 506
rect 344 496 346 501
rect 261 474 267 476
rect 261 472 263 474
rect 265 472 267 474
rect 275 479 277 482
rect 285 479 287 482
rect 305 479 307 482
rect 312 479 314 482
rect 323 479 325 488
rect 357 495 359 500
rect 364 495 366 500
rect 384 496 386 501
rect 397 495 399 500
rect 404 495 406 500
rect 435 499 437 504
rect 475 502 477 506
rect 482 502 484 506
rect 493 502 495 506
rect 445 496 447 501
rect 455 496 457 501
rect 425 486 427 489
rect 425 484 431 486
rect 425 482 427 484
rect 429 482 431 484
rect 344 479 346 482
rect 357 479 359 482
rect 275 477 281 479
rect 275 475 277 477
rect 279 475 281 477
rect 275 473 281 475
rect 285 477 307 479
rect 285 475 296 477
rect 298 475 303 477
rect 305 475 307 477
rect 285 473 307 475
rect 311 477 317 479
rect 311 475 313 477
rect 315 475 317 477
rect 311 473 317 475
rect 321 477 327 479
rect 321 475 323 477
rect 325 475 327 477
rect 321 473 327 475
rect 344 477 350 479
rect 344 475 346 477
rect 348 475 350 477
rect 344 473 350 475
rect 354 477 360 479
rect 354 475 356 477
rect 358 475 360 477
rect 354 473 360 475
rect 261 470 270 472
rect 278 470 280 473
rect 285 470 287 473
rect 303 470 305 473
rect 313 470 315 473
rect 323 470 325 473
rect 344 470 346 473
rect 268 467 270 470
rect 214 449 216 454
rect 78 438 80 442
rect 88 438 90 442
rect 98 438 100 442
rect 118 438 120 442
rect 128 438 130 442
rect 138 438 140 442
rect 159 438 161 442
rect 169 438 171 442
rect 179 438 181 442
rect 197 440 199 445
rect 204 440 206 445
rect 268 449 270 454
rect 227 438 229 442
rect 255 438 257 442
rect 278 440 280 445
rect 285 440 287 445
rect 354 461 356 473
rect 364 471 366 482
rect 384 479 386 482
rect 397 479 399 482
rect 384 477 390 479
rect 384 475 386 477
rect 388 475 390 477
rect 384 473 390 475
rect 394 477 400 479
rect 394 475 396 477
rect 398 475 400 477
rect 394 473 400 475
rect 364 469 370 471
rect 384 470 386 473
rect 364 467 366 469
rect 368 467 370 469
rect 364 465 370 467
rect 364 461 366 465
rect 394 461 396 473
rect 404 471 406 482
rect 425 480 431 482
rect 404 469 410 471
rect 404 467 406 469
rect 408 467 410 469
rect 425 467 427 480
rect 435 476 437 489
rect 514 496 516 501
rect 431 474 437 476
rect 431 472 433 474
rect 435 472 437 474
rect 445 479 447 482
rect 455 479 457 482
rect 475 479 477 482
rect 482 479 484 482
rect 493 479 495 488
rect 527 495 529 500
rect 534 495 536 500
rect 554 496 556 501
rect 675 502 677 506
rect 686 502 688 506
rect 693 502 695 506
rect 567 495 569 500
rect 574 495 576 500
rect 594 495 596 500
rect 601 495 603 500
rect 614 496 616 501
rect 634 495 636 500
rect 641 495 643 500
rect 654 496 656 501
rect 514 479 516 482
rect 527 479 529 482
rect 445 477 451 479
rect 445 475 447 477
rect 449 475 451 477
rect 445 473 451 475
rect 455 477 477 479
rect 455 475 466 477
rect 468 475 473 477
rect 475 475 477 477
rect 455 473 477 475
rect 481 477 487 479
rect 481 475 483 477
rect 485 475 487 477
rect 481 473 487 475
rect 491 477 497 479
rect 491 475 493 477
rect 495 475 497 477
rect 491 473 497 475
rect 514 477 520 479
rect 514 475 516 477
rect 518 475 520 477
rect 514 473 520 475
rect 524 477 530 479
rect 524 475 526 477
rect 528 475 530 477
rect 524 473 530 475
rect 431 470 440 472
rect 448 470 450 473
rect 455 470 457 473
rect 473 470 475 473
rect 483 470 485 473
rect 493 470 495 473
rect 514 470 516 473
rect 438 467 440 470
rect 404 465 410 467
rect 404 461 406 465
rect 438 449 440 454
rect 303 438 305 442
rect 313 438 315 442
rect 323 438 325 442
rect 344 438 346 442
rect 354 438 356 442
rect 364 438 366 442
rect 384 438 386 442
rect 394 438 396 442
rect 404 438 406 442
rect 425 438 427 442
rect 448 440 450 445
rect 455 440 457 445
rect 524 461 526 473
rect 534 471 536 482
rect 554 479 556 482
rect 567 479 569 482
rect 554 477 560 479
rect 554 475 556 477
rect 558 475 560 477
rect 554 473 560 475
rect 564 477 570 479
rect 564 475 566 477
rect 568 475 570 477
rect 564 473 570 475
rect 534 469 540 471
rect 554 470 556 473
rect 534 467 536 469
rect 538 467 540 469
rect 534 465 540 467
rect 534 461 536 465
rect 564 461 566 473
rect 574 471 576 482
rect 594 471 596 482
rect 601 479 603 482
rect 614 479 616 482
rect 600 477 606 479
rect 600 475 602 477
rect 604 475 606 477
rect 600 473 606 475
rect 610 477 616 479
rect 610 475 612 477
rect 614 475 616 477
rect 610 473 616 475
rect 574 469 580 471
rect 574 467 576 469
rect 578 467 580 469
rect 574 465 580 467
rect 590 469 596 471
rect 590 467 592 469
rect 594 467 596 469
rect 590 465 596 467
rect 574 461 576 465
rect 594 461 596 465
rect 604 461 606 473
rect 614 470 616 473
rect 634 471 636 482
rect 641 479 643 482
rect 654 479 656 482
rect 675 479 677 488
rect 713 496 715 501
rect 723 496 725 501
rect 733 499 735 504
rect 743 502 745 506
rect 686 479 688 482
rect 693 479 695 482
rect 713 479 715 482
rect 723 479 725 482
rect 640 477 646 479
rect 640 475 642 477
rect 644 475 646 477
rect 640 473 646 475
rect 650 477 656 479
rect 650 475 652 477
rect 654 475 656 477
rect 650 473 656 475
rect 673 477 679 479
rect 673 475 675 477
rect 677 475 679 477
rect 673 473 679 475
rect 683 477 689 479
rect 683 475 685 477
rect 687 475 689 477
rect 683 473 689 475
rect 693 477 715 479
rect 693 475 695 477
rect 697 475 702 477
rect 704 475 715 477
rect 693 473 715 475
rect 719 477 725 479
rect 719 475 721 477
rect 723 475 725 477
rect 719 473 725 475
rect 733 476 735 489
rect 743 486 745 489
rect 739 484 745 486
rect 739 482 741 484
rect 743 482 745 484
rect 739 480 745 482
rect 733 474 739 476
rect 630 469 636 471
rect 630 467 632 469
rect 634 467 636 469
rect 630 465 636 467
rect 634 461 636 465
rect 644 461 646 473
rect 654 470 656 473
rect 675 470 677 473
rect 685 470 687 473
rect 695 470 697 473
rect 713 470 715 473
rect 720 470 722 473
rect 733 472 735 474
rect 737 472 739 474
rect 730 470 739 472
rect 730 467 732 470
rect 743 467 745 480
rect 730 449 732 454
rect 473 438 475 442
rect 483 438 485 442
rect 493 438 495 442
rect 514 438 516 442
rect 524 438 526 442
rect 534 438 536 442
rect 554 438 556 442
rect 564 438 566 442
rect 574 438 576 442
rect 594 438 596 442
rect 604 438 606 442
rect 614 438 616 442
rect 634 438 636 442
rect 644 438 646 442
rect 654 438 656 442
rect 675 438 677 442
rect 685 438 687 442
rect 695 438 697 442
rect 713 440 715 445
rect 720 440 722 445
rect 743 438 745 442
rect 78 430 80 434
rect 91 430 93 434
rect 98 430 100 434
rect 119 430 121 434
rect 129 430 131 434
rect 139 430 141 434
rect 157 427 159 432
rect 164 427 166 432
rect 187 430 189 434
rect 220 430 222 434
rect 230 430 232 434
rect 240 430 242 434
rect 174 418 176 423
rect 174 402 176 405
rect 78 399 80 402
rect 91 399 93 402
rect 98 399 100 402
rect 119 399 121 402
rect 129 399 131 402
rect 139 399 141 402
rect 157 399 159 402
rect 164 399 166 402
rect 174 400 183 402
rect 78 397 84 399
rect 78 395 80 397
rect 82 395 84 397
rect 78 393 84 395
rect 88 397 94 399
rect 88 395 90 397
rect 92 395 94 397
rect 88 393 94 395
rect 98 397 107 399
rect 98 395 103 397
rect 105 395 107 397
rect 98 393 107 395
rect 117 397 123 399
rect 117 395 119 397
rect 121 395 123 397
rect 117 393 123 395
rect 127 397 133 399
rect 127 395 129 397
rect 131 395 133 397
rect 127 393 133 395
rect 137 397 159 399
rect 137 395 139 397
rect 141 395 146 397
rect 148 395 159 397
rect 137 393 159 395
rect 163 397 169 399
rect 163 395 165 397
rect 167 395 169 397
rect 163 393 169 395
rect 78 390 80 393
rect 88 385 90 393
rect 98 387 100 393
rect 119 384 121 393
rect 130 390 132 393
rect 137 390 139 393
rect 157 390 159 393
rect 167 390 169 393
rect 177 398 179 400
rect 181 398 183 400
rect 177 396 183 398
rect 78 371 80 376
rect 88 372 90 377
rect 98 375 100 379
rect 177 383 179 396
rect 187 392 189 405
rect 258 427 260 432
rect 265 427 267 432
rect 288 430 290 434
rect 322 430 324 434
rect 332 430 334 434
rect 342 430 344 434
rect 275 418 277 423
rect 275 402 277 405
rect 220 399 222 402
rect 230 399 232 402
rect 240 399 242 402
rect 258 399 260 402
rect 265 399 267 402
rect 275 400 284 402
rect 218 397 224 399
rect 218 395 220 397
rect 222 395 224 397
rect 218 393 224 395
rect 228 397 234 399
rect 228 395 230 397
rect 232 395 234 397
rect 228 393 234 395
rect 238 397 260 399
rect 238 395 240 397
rect 242 395 247 397
rect 249 395 260 397
rect 238 393 260 395
rect 264 397 270 399
rect 264 395 266 397
rect 268 395 270 397
rect 264 393 270 395
rect 183 390 189 392
rect 183 388 185 390
rect 187 388 189 390
rect 183 386 189 388
rect 187 383 189 386
rect 220 384 222 393
rect 231 390 233 393
rect 238 390 240 393
rect 258 390 260 393
rect 268 390 270 393
rect 278 398 280 400
rect 282 398 284 400
rect 278 396 284 398
rect 157 371 159 376
rect 167 371 169 376
rect 119 366 121 370
rect 130 366 132 370
rect 137 366 139 370
rect 177 368 179 373
rect 278 383 280 396
rect 288 392 290 405
rect 360 427 362 432
rect 367 427 369 432
rect 390 430 392 434
rect 422 430 424 434
rect 377 418 379 423
rect 377 402 379 405
rect 322 399 324 402
rect 332 399 334 402
rect 342 399 344 402
rect 360 399 362 402
rect 367 399 369 402
rect 377 400 386 402
rect 320 397 326 399
rect 320 395 322 397
rect 324 395 326 397
rect 320 393 326 395
rect 330 397 336 399
rect 330 395 332 397
rect 334 395 336 397
rect 330 393 336 395
rect 340 397 362 399
rect 340 395 342 397
rect 344 395 349 397
rect 351 395 362 397
rect 340 393 362 395
rect 366 397 372 399
rect 366 395 368 397
rect 370 395 372 397
rect 366 393 372 395
rect 284 390 290 392
rect 284 388 286 390
rect 288 388 290 390
rect 284 386 290 388
rect 288 383 290 386
rect 322 384 324 393
rect 333 390 335 393
rect 340 390 342 393
rect 360 390 362 393
rect 370 390 372 393
rect 380 398 382 400
rect 384 398 386 400
rect 380 396 386 398
rect 258 371 260 376
rect 268 371 270 376
rect 187 366 189 370
rect 220 366 222 370
rect 231 366 233 370
rect 238 366 240 370
rect 278 368 280 373
rect 380 383 382 396
rect 390 392 392 405
rect 435 430 437 434
rect 442 430 444 434
rect 475 430 477 434
rect 485 430 487 434
rect 495 430 497 434
rect 513 427 515 432
rect 520 427 522 432
rect 543 430 545 434
rect 576 430 578 434
rect 586 430 588 434
rect 596 430 598 434
rect 530 418 532 423
rect 530 402 532 405
rect 386 390 392 392
rect 422 399 424 402
rect 435 399 437 402
rect 442 399 444 402
rect 475 399 477 402
rect 485 399 487 402
rect 495 399 497 402
rect 513 399 515 402
rect 520 399 522 402
rect 530 400 539 402
rect 422 397 428 399
rect 422 395 424 397
rect 426 395 428 397
rect 422 393 428 395
rect 432 397 438 399
rect 432 395 434 397
rect 436 395 438 397
rect 432 393 438 395
rect 442 397 451 399
rect 442 395 447 397
rect 449 395 451 397
rect 442 393 451 395
rect 473 397 479 399
rect 473 395 475 397
rect 477 395 479 397
rect 473 393 479 395
rect 483 397 489 399
rect 483 395 485 397
rect 487 395 489 397
rect 483 393 489 395
rect 493 397 515 399
rect 493 395 495 397
rect 497 395 502 397
rect 504 395 515 397
rect 493 393 515 395
rect 519 397 525 399
rect 519 395 521 397
rect 523 395 525 397
rect 519 393 525 395
rect 422 390 424 393
rect 386 388 388 390
rect 390 388 392 390
rect 386 386 392 388
rect 390 383 392 386
rect 360 371 362 376
rect 370 371 372 376
rect 288 366 290 370
rect 322 366 324 370
rect 333 366 335 370
rect 340 366 342 370
rect 380 368 382 373
rect 432 385 434 393
rect 442 387 444 393
rect 475 384 477 393
rect 486 390 488 393
rect 493 390 495 393
rect 513 390 515 393
rect 523 390 525 393
rect 533 398 535 400
rect 537 398 539 400
rect 533 396 539 398
rect 422 371 424 376
rect 432 372 434 377
rect 442 375 444 379
rect 390 366 392 370
rect 533 383 535 396
rect 543 392 545 405
rect 614 427 616 432
rect 621 427 623 432
rect 644 430 646 434
rect 675 430 677 434
rect 685 430 687 434
rect 695 430 697 434
rect 631 418 633 423
rect 631 402 633 405
rect 576 399 578 402
rect 586 399 588 402
rect 596 399 598 402
rect 614 399 616 402
rect 621 399 623 402
rect 631 400 640 402
rect 574 397 580 399
rect 574 395 576 397
rect 578 395 580 397
rect 574 393 580 395
rect 584 397 590 399
rect 584 395 586 397
rect 588 395 590 397
rect 584 393 590 395
rect 594 397 616 399
rect 594 395 596 397
rect 598 395 603 397
rect 605 395 616 397
rect 594 393 616 395
rect 620 397 626 399
rect 620 395 622 397
rect 624 395 626 397
rect 620 393 626 395
rect 539 390 545 392
rect 539 388 541 390
rect 543 388 545 390
rect 539 386 545 388
rect 543 383 545 386
rect 576 384 578 393
rect 587 390 589 393
rect 594 390 596 393
rect 614 390 616 393
rect 624 390 626 393
rect 634 398 636 400
rect 638 398 640 400
rect 634 396 640 398
rect 513 371 515 376
rect 523 371 525 376
rect 475 366 477 370
rect 486 366 488 370
rect 493 366 495 370
rect 533 368 535 373
rect 634 383 636 396
rect 644 392 646 405
rect 713 427 715 432
rect 720 427 722 432
rect 743 430 745 434
rect 730 418 732 423
rect 730 402 732 405
rect 675 399 677 402
rect 685 399 687 402
rect 695 399 697 402
rect 713 399 715 402
rect 720 399 722 402
rect 730 400 739 402
rect 673 397 679 399
rect 673 395 675 397
rect 677 395 679 397
rect 673 393 679 395
rect 683 397 689 399
rect 683 395 685 397
rect 687 395 689 397
rect 683 393 689 395
rect 693 397 715 399
rect 693 395 695 397
rect 697 395 702 397
rect 704 395 715 397
rect 693 393 715 395
rect 719 397 725 399
rect 719 395 721 397
rect 723 395 725 397
rect 719 393 725 395
rect 640 390 646 392
rect 640 388 642 390
rect 644 388 646 390
rect 640 386 646 388
rect 644 383 646 386
rect 675 384 677 393
rect 686 390 688 393
rect 693 390 695 393
rect 713 390 715 393
rect 723 390 725 393
rect 733 398 735 400
rect 737 398 739 400
rect 733 396 739 398
rect 614 371 616 376
rect 624 371 626 376
rect 543 366 545 370
rect 576 366 578 370
rect 587 366 589 370
rect 594 366 596 370
rect 634 368 636 373
rect 733 383 735 396
rect 743 392 745 405
rect 739 390 745 392
rect 739 388 741 390
rect 743 388 745 390
rect 739 386 745 388
rect 743 383 745 386
rect 713 371 715 376
rect 723 371 725 376
rect 644 366 646 370
rect 675 366 677 370
rect 686 366 688 370
rect 693 366 695 370
rect 733 368 735 373
rect 743 366 745 370
rect 80 358 82 362
rect 91 358 93 362
rect 98 358 100 362
rect 80 335 82 344
rect 118 352 120 357
rect 128 352 130 357
rect 138 355 140 360
rect 148 358 150 362
rect 221 358 223 362
rect 232 358 234 362
rect 239 358 241 362
rect 168 352 170 357
rect 91 335 93 338
rect 98 335 100 338
rect 118 335 120 338
rect 128 335 130 338
rect 78 333 84 335
rect 78 331 80 333
rect 82 331 84 333
rect 78 329 84 331
rect 88 333 94 335
rect 88 331 90 333
rect 92 331 94 333
rect 88 329 94 331
rect 98 333 120 335
rect 98 331 100 333
rect 102 331 107 333
rect 109 331 120 333
rect 98 329 120 331
rect 124 333 130 335
rect 124 331 126 333
rect 128 331 130 333
rect 124 329 130 331
rect 138 332 140 345
rect 148 342 150 345
rect 144 340 150 342
rect 144 338 146 340
rect 148 338 150 340
rect 178 351 180 356
rect 188 349 190 353
rect 144 336 150 338
rect 138 330 144 332
rect 80 326 82 329
rect 90 326 92 329
rect 100 326 102 329
rect 118 326 120 329
rect 125 326 127 329
rect 138 328 140 330
rect 142 328 144 330
rect 135 326 144 328
rect 135 323 137 326
rect 148 323 150 336
rect 168 335 170 338
rect 178 335 180 343
rect 188 335 190 341
rect 221 335 223 344
rect 259 352 261 357
rect 269 352 271 357
rect 279 355 281 360
rect 289 358 291 362
rect 321 358 323 362
rect 331 355 333 360
rect 371 358 373 362
rect 378 358 380 362
rect 389 358 391 362
rect 341 352 343 357
rect 351 352 353 357
rect 232 335 234 338
rect 239 335 241 338
rect 259 335 261 338
rect 269 335 271 338
rect 168 333 174 335
rect 168 331 170 333
rect 172 331 174 333
rect 168 329 174 331
rect 178 333 184 335
rect 178 331 180 333
rect 182 331 184 333
rect 178 329 184 331
rect 188 333 197 335
rect 188 331 193 333
rect 195 331 197 333
rect 188 329 197 331
rect 219 333 225 335
rect 219 331 221 333
rect 223 331 225 333
rect 219 329 225 331
rect 229 333 235 335
rect 229 331 231 333
rect 233 331 235 333
rect 229 329 235 331
rect 239 333 261 335
rect 239 331 241 333
rect 243 331 248 333
rect 250 331 261 333
rect 239 329 261 331
rect 265 333 271 335
rect 265 331 267 333
rect 269 331 271 333
rect 265 329 271 331
rect 279 332 281 345
rect 289 342 291 345
rect 285 340 291 342
rect 285 338 287 340
rect 289 338 291 340
rect 285 336 291 338
rect 279 330 285 332
rect 168 326 170 329
rect 181 326 183 329
rect 188 326 190 329
rect 221 326 223 329
rect 231 326 233 329
rect 241 326 243 329
rect 259 326 261 329
rect 266 326 268 329
rect 279 328 281 330
rect 283 328 285 330
rect 276 326 285 328
rect 135 305 137 310
rect 80 294 82 298
rect 90 294 92 298
rect 100 294 102 298
rect 118 296 120 301
rect 125 296 127 301
rect 148 294 150 298
rect 168 294 170 298
rect 276 323 278 326
rect 289 323 291 336
rect 321 342 323 345
rect 321 340 327 342
rect 321 338 323 340
rect 325 338 327 340
rect 321 336 327 338
rect 321 323 323 336
rect 331 332 333 345
rect 475 358 477 362
rect 486 358 488 362
rect 493 358 495 362
rect 422 352 424 357
rect 327 330 333 332
rect 327 328 329 330
rect 331 328 333 330
rect 341 335 343 338
rect 351 335 353 338
rect 371 335 373 338
rect 378 335 380 338
rect 389 335 391 344
rect 432 351 434 356
rect 442 349 444 353
rect 422 335 424 338
rect 432 335 434 343
rect 442 335 444 341
rect 475 335 477 344
rect 513 352 515 357
rect 523 352 525 357
rect 533 355 535 360
rect 543 358 545 362
rect 576 358 578 362
rect 587 358 589 362
rect 594 358 596 362
rect 486 335 488 338
rect 493 335 495 338
rect 513 335 515 338
rect 523 335 525 338
rect 341 333 347 335
rect 341 331 343 333
rect 345 331 347 333
rect 341 329 347 331
rect 351 333 373 335
rect 351 331 362 333
rect 364 331 369 333
rect 371 331 373 333
rect 351 329 373 331
rect 377 333 383 335
rect 377 331 379 333
rect 381 331 383 333
rect 377 329 383 331
rect 387 333 393 335
rect 387 331 389 333
rect 391 331 393 333
rect 387 329 393 331
rect 422 333 428 335
rect 422 331 424 333
rect 426 331 428 333
rect 422 329 428 331
rect 432 333 438 335
rect 432 331 434 333
rect 436 331 438 333
rect 432 329 438 331
rect 442 333 451 335
rect 442 331 447 333
rect 449 331 451 333
rect 442 329 451 331
rect 473 333 479 335
rect 473 331 475 333
rect 477 331 479 333
rect 473 329 479 331
rect 483 333 489 335
rect 483 331 485 333
rect 487 331 489 333
rect 483 329 489 331
rect 493 333 515 335
rect 493 331 495 333
rect 497 331 502 333
rect 504 331 515 333
rect 493 329 515 331
rect 519 333 525 335
rect 519 331 521 333
rect 523 331 525 333
rect 519 329 525 331
rect 533 332 535 345
rect 543 342 545 345
rect 539 340 545 342
rect 539 338 541 340
rect 543 338 545 340
rect 539 336 545 338
rect 533 330 539 332
rect 327 326 336 328
rect 344 326 346 329
rect 351 326 353 329
rect 369 326 371 329
rect 379 326 381 329
rect 389 326 391 329
rect 422 326 424 329
rect 435 326 437 329
rect 442 326 444 329
rect 475 326 477 329
rect 485 326 487 329
rect 495 326 497 329
rect 513 326 515 329
rect 520 326 522 329
rect 533 328 535 330
rect 537 328 539 330
rect 530 326 539 328
rect 334 323 336 326
rect 276 305 278 310
rect 181 294 183 298
rect 188 294 190 298
rect 221 294 223 298
rect 231 294 233 298
rect 241 294 243 298
rect 259 296 261 301
rect 266 296 268 301
rect 334 305 336 310
rect 289 294 291 298
rect 321 294 323 298
rect 344 296 346 301
rect 351 296 353 301
rect 369 294 371 298
rect 379 294 381 298
rect 389 294 391 298
rect 422 294 424 298
rect 530 323 532 326
rect 543 323 545 336
rect 576 335 578 344
rect 614 352 616 357
rect 624 352 626 357
rect 634 355 636 360
rect 644 358 646 362
rect 675 358 677 362
rect 686 358 688 362
rect 693 358 695 362
rect 587 335 589 338
rect 594 335 596 338
rect 614 335 616 338
rect 624 335 626 338
rect 574 333 580 335
rect 574 331 576 333
rect 578 331 580 333
rect 574 329 580 331
rect 584 333 590 335
rect 584 331 586 333
rect 588 331 590 333
rect 584 329 590 331
rect 594 333 616 335
rect 594 331 596 333
rect 598 331 603 333
rect 605 331 616 333
rect 594 329 616 331
rect 620 333 626 335
rect 620 331 622 333
rect 624 331 626 333
rect 620 329 626 331
rect 634 332 636 345
rect 644 342 646 345
rect 640 340 646 342
rect 640 338 642 340
rect 644 338 646 340
rect 640 336 646 338
rect 634 330 640 332
rect 576 326 578 329
rect 586 326 588 329
rect 596 326 598 329
rect 614 326 616 329
rect 621 326 623 329
rect 634 328 636 330
rect 638 328 640 330
rect 631 326 640 328
rect 530 305 532 310
rect 435 294 437 298
rect 442 294 444 298
rect 475 294 477 298
rect 485 294 487 298
rect 495 294 497 298
rect 513 296 515 301
rect 520 296 522 301
rect 631 323 633 326
rect 644 323 646 336
rect 675 335 677 344
rect 713 352 715 357
rect 723 352 725 357
rect 733 355 735 360
rect 743 358 745 362
rect 686 335 688 338
rect 693 335 695 338
rect 713 335 715 338
rect 723 335 725 338
rect 673 333 679 335
rect 673 331 675 333
rect 677 331 679 333
rect 673 329 679 331
rect 683 333 689 335
rect 683 331 685 333
rect 687 331 689 333
rect 683 329 689 331
rect 693 333 715 335
rect 693 331 695 333
rect 697 331 702 333
rect 704 331 715 333
rect 693 329 715 331
rect 719 333 725 335
rect 719 331 721 333
rect 723 331 725 333
rect 719 329 725 331
rect 733 332 735 345
rect 743 342 745 345
rect 739 340 745 342
rect 739 338 741 340
rect 743 338 745 340
rect 739 336 745 338
rect 733 330 739 332
rect 675 326 677 329
rect 685 326 687 329
rect 695 326 697 329
rect 713 326 715 329
rect 720 326 722 329
rect 733 328 735 330
rect 737 328 739 330
rect 730 326 739 328
rect 631 305 633 310
rect 543 294 545 298
rect 576 294 578 298
rect 586 294 588 298
rect 596 294 598 298
rect 614 296 616 301
rect 621 296 623 301
rect 730 323 732 326
rect 743 323 745 336
rect 730 305 732 310
rect 644 294 646 298
rect 675 294 677 298
rect 685 294 687 298
rect 695 294 697 298
rect 713 296 715 301
rect 720 296 722 301
rect 743 294 745 298
rect 78 286 80 290
rect 91 286 93 290
rect 98 286 100 290
rect 119 286 121 290
rect 129 286 131 290
rect 139 286 141 290
rect 157 283 159 288
rect 164 283 166 288
rect 187 286 189 290
rect 220 286 222 290
rect 230 286 232 290
rect 240 286 242 290
rect 174 274 176 279
rect 174 258 176 261
rect 78 255 80 258
rect 91 255 93 258
rect 98 255 100 258
rect 119 255 121 258
rect 129 255 131 258
rect 139 255 141 258
rect 157 255 159 258
rect 164 255 166 258
rect 174 256 183 258
rect 78 253 84 255
rect 78 251 80 253
rect 82 251 84 253
rect 78 249 84 251
rect 88 253 94 255
rect 88 251 90 253
rect 92 251 94 253
rect 88 249 94 251
rect 98 253 107 255
rect 98 251 103 253
rect 105 251 107 253
rect 98 249 107 251
rect 117 253 123 255
rect 117 251 119 253
rect 121 251 123 253
rect 117 249 123 251
rect 127 253 133 255
rect 127 251 129 253
rect 131 251 133 253
rect 127 249 133 251
rect 137 253 159 255
rect 137 251 139 253
rect 141 251 146 253
rect 148 251 159 253
rect 137 249 159 251
rect 163 253 169 255
rect 163 251 165 253
rect 167 251 169 253
rect 163 249 169 251
rect 78 246 80 249
rect 88 241 90 249
rect 98 243 100 249
rect 119 240 121 249
rect 130 246 132 249
rect 137 246 139 249
rect 157 246 159 249
rect 167 246 169 249
rect 177 254 179 256
rect 181 254 183 256
rect 177 252 183 254
rect 78 227 80 232
rect 88 228 90 233
rect 98 231 100 235
rect 177 239 179 252
rect 187 248 189 261
rect 258 283 260 288
rect 265 283 267 288
rect 288 286 290 290
rect 321 286 323 290
rect 331 286 333 290
rect 341 286 343 290
rect 275 274 277 279
rect 275 258 277 261
rect 220 255 222 258
rect 230 255 232 258
rect 240 255 242 258
rect 258 255 260 258
rect 265 255 267 258
rect 275 256 284 258
rect 218 253 224 255
rect 218 251 220 253
rect 222 251 224 253
rect 218 249 224 251
rect 228 253 234 255
rect 228 251 230 253
rect 232 251 234 253
rect 228 249 234 251
rect 238 253 260 255
rect 238 251 240 253
rect 242 251 247 253
rect 249 251 260 253
rect 238 249 260 251
rect 264 253 270 255
rect 264 251 266 253
rect 268 251 270 253
rect 264 249 270 251
rect 183 246 189 248
rect 183 244 185 246
rect 187 244 189 246
rect 183 242 189 244
rect 187 239 189 242
rect 220 240 222 249
rect 231 246 233 249
rect 238 246 240 249
rect 258 246 260 249
rect 268 246 270 249
rect 278 254 280 256
rect 282 254 284 256
rect 278 252 284 254
rect 157 227 159 232
rect 167 227 169 232
rect 119 222 121 226
rect 130 222 132 226
rect 137 222 139 226
rect 177 224 179 229
rect 278 239 280 252
rect 288 248 290 261
rect 359 283 361 288
rect 366 283 368 288
rect 389 286 391 290
rect 421 286 423 290
rect 376 274 378 279
rect 376 258 378 261
rect 321 255 323 258
rect 331 255 333 258
rect 341 255 343 258
rect 359 255 361 258
rect 366 255 368 258
rect 376 256 385 258
rect 319 253 325 255
rect 319 251 321 253
rect 323 251 325 253
rect 319 249 325 251
rect 329 253 335 255
rect 329 251 331 253
rect 333 251 335 253
rect 329 249 335 251
rect 339 253 361 255
rect 339 251 341 253
rect 343 251 348 253
rect 350 251 361 253
rect 339 249 361 251
rect 365 253 371 255
rect 365 251 367 253
rect 369 251 371 253
rect 365 249 371 251
rect 284 246 290 248
rect 284 244 286 246
rect 288 244 290 246
rect 284 242 290 244
rect 288 239 290 242
rect 321 240 323 249
rect 332 246 334 249
rect 339 246 341 249
rect 359 246 361 249
rect 369 246 371 249
rect 379 254 381 256
rect 383 254 385 256
rect 379 252 385 254
rect 258 227 260 232
rect 268 227 270 232
rect 187 222 189 226
rect 220 222 222 226
rect 231 222 233 226
rect 238 222 240 226
rect 278 224 280 229
rect 379 239 381 252
rect 389 248 391 261
rect 434 286 436 290
rect 441 286 443 290
rect 474 286 476 290
rect 484 286 486 290
rect 494 286 496 290
rect 512 283 514 288
rect 519 283 521 288
rect 542 286 544 290
rect 575 286 577 290
rect 585 286 587 290
rect 595 286 597 290
rect 529 274 531 279
rect 529 258 531 261
rect 385 246 391 248
rect 421 255 423 258
rect 434 255 436 258
rect 441 255 443 258
rect 474 255 476 258
rect 484 255 486 258
rect 494 255 496 258
rect 512 255 514 258
rect 519 255 521 258
rect 529 256 538 258
rect 421 253 427 255
rect 421 251 423 253
rect 425 251 427 253
rect 421 249 427 251
rect 431 253 437 255
rect 431 251 433 253
rect 435 251 437 253
rect 431 249 437 251
rect 441 253 450 255
rect 441 251 446 253
rect 448 251 450 253
rect 441 249 450 251
rect 472 253 478 255
rect 472 251 474 253
rect 476 251 478 253
rect 472 249 478 251
rect 482 253 488 255
rect 482 251 484 253
rect 486 251 488 253
rect 482 249 488 251
rect 492 253 514 255
rect 492 251 494 253
rect 496 251 501 253
rect 503 251 514 253
rect 492 249 514 251
rect 518 253 524 255
rect 518 251 520 253
rect 522 251 524 253
rect 518 249 524 251
rect 421 246 423 249
rect 385 244 387 246
rect 389 244 391 246
rect 385 242 391 244
rect 389 239 391 242
rect 359 227 361 232
rect 369 227 371 232
rect 288 222 290 226
rect 321 222 323 226
rect 332 222 334 226
rect 339 222 341 226
rect 379 224 381 229
rect 431 241 433 249
rect 441 243 443 249
rect 474 240 476 249
rect 485 246 487 249
rect 492 246 494 249
rect 512 246 514 249
rect 522 246 524 249
rect 532 254 534 256
rect 536 254 538 256
rect 532 252 538 254
rect 421 227 423 232
rect 431 228 433 233
rect 441 231 443 235
rect 389 222 391 226
rect 532 239 534 252
rect 542 248 544 261
rect 613 283 615 288
rect 620 283 622 288
rect 643 286 645 290
rect 674 286 676 290
rect 684 286 686 290
rect 694 286 696 290
rect 630 274 632 279
rect 630 258 632 261
rect 575 255 577 258
rect 585 255 587 258
rect 595 255 597 258
rect 613 255 615 258
rect 620 255 622 258
rect 630 256 639 258
rect 573 253 579 255
rect 573 251 575 253
rect 577 251 579 253
rect 573 249 579 251
rect 583 253 589 255
rect 583 251 585 253
rect 587 251 589 253
rect 583 249 589 251
rect 593 253 615 255
rect 593 251 595 253
rect 597 251 602 253
rect 604 251 615 253
rect 593 249 615 251
rect 619 253 625 255
rect 619 251 621 253
rect 623 251 625 253
rect 619 249 625 251
rect 538 246 544 248
rect 538 244 540 246
rect 542 244 544 246
rect 538 242 544 244
rect 542 239 544 242
rect 575 240 577 249
rect 586 246 588 249
rect 593 246 595 249
rect 613 246 615 249
rect 623 246 625 249
rect 633 254 635 256
rect 637 254 639 256
rect 633 252 639 254
rect 512 227 514 232
rect 522 227 524 232
rect 474 222 476 226
rect 485 222 487 226
rect 492 222 494 226
rect 532 224 534 229
rect 633 239 635 252
rect 643 248 645 261
rect 712 283 714 288
rect 719 283 721 288
rect 742 286 744 290
rect 729 274 731 279
rect 729 258 731 261
rect 674 255 676 258
rect 684 255 686 258
rect 694 255 696 258
rect 712 255 714 258
rect 719 255 721 258
rect 729 256 738 258
rect 672 253 678 255
rect 672 251 674 253
rect 676 251 678 253
rect 672 249 678 251
rect 682 253 688 255
rect 682 251 684 253
rect 686 251 688 253
rect 682 249 688 251
rect 692 253 714 255
rect 692 251 694 253
rect 696 251 701 253
rect 703 251 714 253
rect 692 249 714 251
rect 718 253 724 255
rect 718 251 720 253
rect 722 251 724 253
rect 718 249 724 251
rect 639 246 645 248
rect 639 244 641 246
rect 643 244 645 246
rect 639 242 645 244
rect 643 239 645 242
rect 674 240 676 249
rect 685 246 687 249
rect 692 246 694 249
rect 712 246 714 249
rect 722 246 724 249
rect 732 254 734 256
rect 736 254 738 256
rect 732 252 738 254
rect 613 227 615 232
rect 623 227 625 232
rect 542 222 544 226
rect 575 222 577 226
rect 586 222 588 226
rect 593 222 595 226
rect 633 224 635 229
rect 732 239 734 252
rect 742 248 744 261
rect 738 246 744 248
rect 738 244 740 246
rect 742 244 744 246
rect 738 242 744 244
rect 742 239 744 242
rect 712 227 714 232
rect 722 227 724 232
rect 643 222 645 226
rect 674 222 676 226
rect 685 222 687 226
rect 692 222 694 226
rect 732 224 734 229
rect 742 222 744 226
<< ndif >>
rect 73 527 78 534
rect 71 525 78 527
rect 71 523 73 525
rect 75 523 78 525
rect 71 521 78 523
rect 80 521 85 534
rect 87 521 98 534
rect 89 520 98 521
rect 100 532 107 534
rect 100 530 103 532
rect 105 530 107 532
rect 100 524 107 530
rect 113 527 118 534
rect 100 522 103 524
rect 105 522 107 524
rect 100 520 107 522
rect 111 525 118 527
rect 111 523 113 525
rect 115 523 118 525
rect 111 521 118 523
rect 120 521 125 534
rect 127 521 138 534
rect 89 515 96 520
rect 129 520 138 521
rect 140 532 147 534
rect 140 530 143 532
rect 145 530 147 532
rect 140 524 147 530
rect 163 528 170 534
rect 140 522 143 524
rect 145 522 147 524
rect 140 520 147 522
rect 152 525 159 528
rect 152 523 154 525
rect 156 523 159 525
rect 152 521 159 523
rect 129 515 136 520
rect 89 513 92 515
rect 94 513 96 515
rect 89 511 96 513
rect 129 513 132 515
rect 134 513 136 515
rect 154 514 159 521
rect 161 518 170 528
rect 161 516 165 518
rect 167 516 170 518
rect 161 514 170 516
rect 172 514 177 534
rect 179 527 184 534
rect 190 532 197 534
rect 190 530 192 532
rect 194 530 197 532
rect 179 525 186 527
rect 179 523 182 525
rect 184 523 186 525
rect 179 521 186 523
rect 190 525 197 530
rect 190 523 192 525
rect 194 523 197 525
rect 179 514 184 521
rect 190 520 197 523
rect 199 532 207 534
rect 199 530 202 532
rect 204 530 207 532
rect 199 520 207 530
rect 209 527 214 534
rect 270 527 275 534
rect 209 524 217 527
rect 209 522 212 524
rect 214 522 217 524
rect 209 520 217 522
rect 212 517 217 520
rect 219 521 227 527
rect 219 519 222 521
rect 224 519 227 521
rect 219 517 227 519
rect 129 511 136 513
rect 222 514 227 517
rect 229 525 236 527
rect 229 523 232 525
rect 234 523 236 525
rect 229 521 236 523
rect 248 525 255 527
rect 248 523 250 525
rect 252 523 255 525
rect 248 521 255 523
rect 229 514 234 521
rect 250 514 255 521
rect 257 521 265 527
rect 257 519 260 521
rect 262 519 265 521
rect 257 517 265 519
rect 267 524 275 527
rect 267 522 270 524
rect 272 522 275 524
rect 267 520 275 522
rect 277 532 285 534
rect 277 530 280 532
rect 282 530 285 532
rect 277 520 285 530
rect 287 532 294 534
rect 287 530 290 532
rect 292 530 294 532
rect 287 525 294 530
rect 300 527 305 534
rect 287 523 290 525
rect 292 523 294 525
rect 287 520 294 523
rect 298 525 305 527
rect 298 523 300 525
rect 302 523 305 525
rect 298 521 305 523
rect 267 517 272 520
rect 257 514 262 517
rect 300 514 305 521
rect 307 514 312 534
rect 314 528 321 534
rect 337 532 344 534
rect 337 530 339 532
rect 341 530 344 532
rect 314 518 323 528
rect 314 516 317 518
rect 319 516 323 518
rect 314 514 323 516
rect 325 525 332 528
rect 325 523 328 525
rect 330 523 332 525
rect 325 521 332 523
rect 337 524 344 530
rect 337 522 339 524
rect 341 522 344 524
rect 325 514 330 521
rect 337 520 344 522
rect 346 521 357 534
rect 359 521 364 534
rect 366 527 371 534
rect 377 532 384 534
rect 377 530 379 532
rect 381 530 384 532
rect 366 525 373 527
rect 366 523 369 525
rect 371 523 373 525
rect 366 521 373 523
rect 377 524 384 530
rect 377 522 379 524
rect 381 522 384 524
rect 346 520 355 521
rect 348 515 355 520
rect 377 520 384 522
rect 386 521 397 534
rect 399 521 404 534
rect 406 527 411 534
rect 440 527 445 534
rect 406 525 413 527
rect 406 523 409 525
rect 411 523 413 525
rect 406 521 413 523
rect 418 525 425 527
rect 418 523 420 525
rect 422 523 425 525
rect 418 521 425 523
rect 386 520 395 521
rect 388 515 395 520
rect 348 513 350 515
rect 352 513 355 515
rect 348 511 355 513
rect 388 513 390 515
rect 392 513 395 515
rect 420 514 425 521
rect 427 521 435 527
rect 427 519 430 521
rect 432 519 435 521
rect 427 517 435 519
rect 437 524 445 527
rect 437 522 440 524
rect 442 522 445 524
rect 437 520 445 522
rect 447 532 455 534
rect 447 530 450 532
rect 452 530 455 532
rect 447 520 455 530
rect 457 532 464 534
rect 457 530 460 532
rect 462 530 464 532
rect 457 525 464 530
rect 470 527 475 534
rect 457 523 460 525
rect 462 523 464 525
rect 457 520 464 523
rect 468 525 475 527
rect 468 523 470 525
rect 472 523 475 525
rect 468 521 475 523
rect 437 517 442 520
rect 427 514 432 517
rect 388 511 395 513
rect 470 514 475 521
rect 477 514 482 534
rect 484 528 491 534
rect 507 532 514 534
rect 507 530 509 532
rect 511 530 514 532
rect 484 518 493 528
rect 484 516 487 518
rect 489 516 493 518
rect 484 514 493 516
rect 495 525 502 528
rect 495 523 498 525
rect 500 523 502 525
rect 495 521 502 523
rect 507 524 514 530
rect 507 522 509 524
rect 511 522 514 524
rect 495 514 500 521
rect 507 520 514 522
rect 516 521 527 534
rect 529 521 534 534
rect 536 527 541 534
rect 547 532 554 534
rect 547 530 549 532
rect 551 530 554 532
rect 536 525 543 527
rect 536 523 539 525
rect 541 523 543 525
rect 536 521 543 523
rect 547 524 554 530
rect 547 522 549 524
rect 551 522 554 524
rect 516 520 525 521
rect 518 515 525 520
rect 547 520 554 522
rect 556 521 567 534
rect 569 521 574 534
rect 576 527 581 534
rect 589 527 594 534
rect 576 525 583 527
rect 576 523 579 525
rect 581 523 583 525
rect 576 521 583 523
rect 587 525 594 527
rect 587 523 589 525
rect 591 523 594 525
rect 587 521 594 523
rect 596 521 601 534
rect 603 521 614 534
rect 556 520 565 521
rect 558 515 565 520
rect 605 520 614 521
rect 616 532 623 534
rect 616 530 619 532
rect 621 530 623 532
rect 616 524 623 530
rect 629 527 634 534
rect 616 522 619 524
rect 621 522 623 524
rect 616 520 623 522
rect 627 525 634 527
rect 627 523 629 525
rect 631 523 634 525
rect 627 521 634 523
rect 636 521 641 534
rect 643 521 654 534
rect 518 513 520 515
rect 522 513 525 515
rect 518 511 525 513
rect 558 513 560 515
rect 562 513 565 515
rect 558 511 565 513
rect 605 515 612 520
rect 645 520 654 521
rect 656 532 663 534
rect 656 530 659 532
rect 661 530 663 532
rect 656 524 663 530
rect 679 528 686 534
rect 656 522 659 524
rect 661 522 663 524
rect 656 520 663 522
rect 668 525 675 528
rect 668 523 670 525
rect 672 523 675 525
rect 668 521 675 523
rect 645 515 652 520
rect 605 513 608 515
rect 610 513 612 515
rect 605 511 612 513
rect 645 513 648 515
rect 650 513 652 515
rect 670 514 675 521
rect 677 518 686 528
rect 677 516 681 518
rect 683 516 686 518
rect 677 514 686 516
rect 688 514 693 534
rect 695 527 700 534
rect 706 532 713 534
rect 706 530 708 532
rect 710 530 713 532
rect 695 525 702 527
rect 695 523 698 525
rect 700 523 702 525
rect 695 521 702 523
rect 706 525 713 530
rect 706 523 708 525
rect 710 523 713 525
rect 695 514 700 521
rect 706 520 713 523
rect 715 532 723 534
rect 715 530 718 532
rect 720 530 723 532
rect 715 520 723 530
rect 725 527 730 534
rect 725 524 733 527
rect 725 522 728 524
rect 730 522 733 524
rect 725 520 733 522
rect 728 517 733 520
rect 735 521 743 527
rect 735 519 738 521
rect 740 519 743 521
rect 735 517 743 519
rect 645 511 652 513
rect 738 514 743 517
rect 745 525 752 527
rect 745 523 748 525
rect 750 523 752 525
rect 745 521 752 523
rect 745 514 750 521
rect 89 503 96 505
rect 89 501 92 503
rect 94 501 96 503
rect 129 503 136 505
rect 129 501 132 503
rect 134 501 136 503
rect 89 496 96 501
rect 89 495 98 496
rect 71 493 78 495
rect 71 491 73 493
rect 75 491 78 493
rect 71 489 78 491
rect 73 482 78 489
rect 80 482 85 495
rect 87 482 98 495
rect 100 494 107 496
rect 129 496 136 501
rect 129 495 138 496
rect 100 492 103 494
rect 105 492 107 494
rect 100 486 107 492
rect 111 493 118 495
rect 111 491 113 493
rect 115 491 118 493
rect 111 489 118 491
rect 100 484 103 486
rect 105 484 107 486
rect 100 482 107 484
rect 113 482 118 489
rect 120 482 125 495
rect 127 482 138 495
rect 140 494 147 496
rect 154 495 159 502
rect 140 492 143 494
rect 145 492 147 494
rect 140 486 147 492
rect 152 493 159 495
rect 152 491 154 493
rect 156 491 159 493
rect 152 488 159 491
rect 161 500 170 502
rect 161 498 165 500
rect 167 498 170 500
rect 161 488 170 498
rect 140 484 143 486
rect 145 484 147 486
rect 140 482 147 484
rect 163 482 170 488
rect 172 482 177 502
rect 179 495 184 502
rect 222 499 227 502
rect 212 496 217 499
rect 179 493 186 495
rect 179 491 182 493
rect 184 491 186 493
rect 179 489 186 491
rect 190 493 197 496
rect 190 491 192 493
rect 194 491 197 493
rect 179 482 184 489
rect 190 486 197 491
rect 190 484 192 486
rect 194 484 197 486
rect 190 482 197 484
rect 199 486 207 496
rect 199 484 202 486
rect 204 484 207 486
rect 199 482 207 484
rect 209 494 217 496
rect 209 492 212 494
rect 214 492 217 494
rect 209 489 217 492
rect 219 497 227 499
rect 219 495 222 497
rect 224 495 227 497
rect 219 489 227 495
rect 229 495 234 502
rect 250 495 255 502
rect 229 493 236 495
rect 229 491 232 493
rect 234 491 236 493
rect 229 489 236 491
rect 248 493 255 495
rect 248 491 250 493
rect 252 491 255 493
rect 248 489 255 491
rect 257 499 262 502
rect 348 503 355 505
rect 257 497 265 499
rect 257 495 260 497
rect 262 495 265 497
rect 257 489 265 495
rect 267 496 272 499
rect 267 494 275 496
rect 267 492 270 494
rect 272 492 275 494
rect 267 489 275 492
rect 209 482 214 489
rect 270 482 275 489
rect 277 486 285 496
rect 277 484 280 486
rect 282 484 285 486
rect 277 482 285 484
rect 287 493 294 496
rect 300 495 305 502
rect 287 491 290 493
rect 292 491 294 493
rect 287 486 294 491
rect 298 493 305 495
rect 298 491 300 493
rect 302 491 305 493
rect 298 489 305 491
rect 287 484 290 486
rect 292 484 294 486
rect 287 482 294 484
rect 300 482 305 489
rect 307 482 312 502
rect 314 500 323 502
rect 314 498 317 500
rect 319 498 323 500
rect 314 488 323 498
rect 325 495 330 502
rect 348 501 350 503
rect 352 501 355 503
rect 388 503 395 505
rect 388 501 390 503
rect 392 501 395 503
rect 348 496 355 501
rect 325 493 332 495
rect 325 491 328 493
rect 330 491 332 493
rect 325 488 332 491
rect 337 494 344 496
rect 337 492 339 494
rect 341 492 344 494
rect 314 482 321 488
rect 337 486 344 492
rect 337 484 339 486
rect 341 484 344 486
rect 337 482 344 484
rect 346 495 355 496
rect 388 496 395 501
rect 346 482 357 495
rect 359 482 364 495
rect 366 493 373 495
rect 366 491 369 493
rect 371 491 373 493
rect 366 489 373 491
rect 377 494 384 496
rect 377 492 379 494
rect 381 492 384 494
rect 366 482 371 489
rect 377 486 384 492
rect 377 484 379 486
rect 381 484 384 486
rect 377 482 384 484
rect 386 495 395 496
rect 420 495 425 502
rect 386 482 397 495
rect 399 482 404 495
rect 406 493 413 495
rect 406 491 409 493
rect 411 491 413 493
rect 406 489 413 491
rect 418 493 425 495
rect 418 491 420 493
rect 422 491 425 493
rect 418 489 425 491
rect 427 499 432 502
rect 518 503 525 505
rect 427 497 435 499
rect 427 495 430 497
rect 432 495 435 497
rect 427 489 435 495
rect 437 496 442 499
rect 437 494 445 496
rect 437 492 440 494
rect 442 492 445 494
rect 437 489 445 492
rect 406 482 411 489
rect 440 482 445 489
rect 447 486 455 496
rect 447 484 450 486
rect 452 484 455 486
rect 447 482 455 484
rect 457 493 464 496
rect 470 495 475 502
rect 457 491 460 493
rect 462 491 464 493
rect 457 486 464 491
rect 468 493 475 495
rect 468 491 470 493
rect 472 491 475 493
rect 468 489 475 491
rect 457 484 460 486
rect 462 484 464 486
rect 457 482 464 484
rect 470 482 475 489
rect 477 482 482 502
rect 484 500 493 502
rect 484 498 487 500
rect 489 498 493 500
rect 484 488 493 498
rect 495 495 500 502
rect 518 501 520 503
rect 522 501 525 503
rect 558 503 565 505
rect 558 501 560 503
rect 562 501 565 503
rect 518 496 525 501
rect 495 493 502 495
rect 495 491 498 493
rect 500 491 502 493
rect 495 488 502 491
rect 507 494 514 496
rect 507 492 509 494
rect 511 492 514 494
rect 484 482 491 488
rect 507 486 514 492
rect 507 484 509 486
rect 511 484 514 486
rect 507 482 514 484
rect 516 495 525 496
rect 558 496 565 501
rect 605 503 612 505
rect 605 501 608 503
rect 610 501 612 503
rect 645 503 652 505
rect 645 501 648 503
rect 650 501 652 503
rect 516 482 527 495
rect 529 482 534 495
rect 536 493 543 495
rect 536 491 539 493
rect 541 491 543 493
rect 536 489 543 491
rect 547 494 554 496
rect 547 492 549 494
rect 551 492 554 494
rect 536 482 541 489
rect 547 486 554 492
rect 547 484 549 486
rect 551 484 554 486
rect 547 482 554 484
rect 556 495 565 496
rect 605 496 612 501
rect 605 495 614 496
rect 556 482 567 495
rect 569 482 574 495
rect 576 493 583 495
rect 576 491 579 493
rect 581 491 583 493
rect 576 489 583 491
rect 587 493 594 495
rect 587 491 589 493
rect 591 491 594 493
rect 587 489 594 491
rect 576 482 581 489
rect 589 482 594 489
rect 596 482 601 495
rect 603 482 614 495
rect 616 494 623 496
rect 645 496 652 501
rect 645 495 654 496
rect 616 492 619 494
rect 621 492 623 494
rect 616 486 623 492
rect 627 493 634 495
rect 627 491 629 493
rect 631 491 634 493
rect 627 489 634 491
rect 616 484 619 486
rect 621 484 623 486
rect 616 482 623 484
rect 629 482 634 489
rect 636 482 641 495
rect 643 482 654 495
rect 656 494 663 496
rect 670 495 675 502
rect 656 492 659 494
rect 661 492 663 494
rect 656 486 663 492
rect 668 493 675 495
rect 668 491 670 493
rect 672 491 675 493
rect 668 488 675 491
rect 677 500 686 502
rect 677 498 681 500
rect 683 498 686 500
rect 677 488 686 498
rect 656 484 659 486
rect 661 484 663 486
rect 656 482 663 484
rect 679 482 686 488
rect 688 482 693 502
rect 695 495 700 502
rect 738 499 743 502
rect 728 496 733 499
rect 695 493 702 495
rect 695 491 698 493
rect 700 491 702 493
rect 695 489 702 491
rect 706 493 713 496
rect 706 491 708 493
rect 710 491 713 493
rect 695 482 700 489
rect 706 486 713 491
rect 706 484 708 486
rect 710 484 713 486
rect 706 482 713 484
rect 715 486 723 496
rect 715 484 718 486
rect 720 484 723 486
rect 715 482 723 484
rect 725 494 733 496
rect 725 492 728 494
rect 730 492 733 494
rect 725 489 733 492
rect 735 497 743 499
rect 735 495 738 497
rect 740 495 743 497
rect 735 489 743 495
rect 745 495 750 502
rect 745 493 752 495
rect 745 491 748 493
rect 750 491 752 493
rect 745 489 752 491
rect 725 482 730 489
rect 71 388 78 390
rect 71 386 73 388
rect 75 386 78 388
rect 71 381 78 386
rect 71 379 73 381
rect 75 379 78 381
rect 71 376 78 379
rect 80 385 85 390
rect 93 385 98 387
rect 80 381 88 385
rect 80 379 83 381
rect 85 379 88 381
rect 80 377 88 379
rect 90 383 98 385
rect 90 381 93 383
rect 95 381 98 383
rect 90 379 98 381
rect 100 383 107 387
rect 123 384 130 390
rect 100 381 103 383
rect 105 381 107 383
rect 100 379 107 381
rect 112 381 119 384
rect 112 379 114 381
rect 116 379 119 381
rect 90 377 95 379
rect 80 376 85 377
rect 112 377 119 379
rect 114 370 119 377
rect 121 374 130 384
rect 121 372 125 374
rect 127 372 130 374
rect 121 370 130 372
rect 132 370 137 390
rect 139 383 144 390
rect 150 388 157 390
rect 150 386 152 388
rect 154 386 157 388
rect 139 381 146 383
rect 139 379 142 381
rect 144 379 146 381
rect 139 377 146 379
rect 150 381 157 386
rect 150 379 152 381
rect 154 379 157 381
rect 139 370 144 377
rect 150 376 157 379
rect 159 388 167 390
rect 159 386 162 388
rect 164 386 167 388
rect 159 376 167 386
rect 169 383 174 390
rect 224 384 231 390
rect 169 380 177 383
rect 169 378 172 380
rect 174 378 177 380
rect 169 376 177 378
rect 172 373 177 376
rect 179 377 187 383
rect 179 375 182 377
rect 184 375 187 377
rect 179 373 187 375
rect 182 370 187 373
rect 189 381 196 383
rect 189 379 192 381
rect 194 379 196 381
rect 189 377 196 379
rect 213 381 220 384
rect 213 379 215 381
rect 217 379 220 381
rect 213 377 220 379
rect 189 370 194 377
rect 215 370 220 377
rect 222 374 231 384
rect 222 372 226 374
rect 228 372 231 374
rect 222 370 231 372
rect 233 370 238 390
rect 240 383 245 390
rect 251 388 258 390
rect 251 386 253 388
rect 255 386 258 388
rect 240 381 247 383
rect 240 379 243 381
rect 245 379 247 381
rect 240 377 247 379
rect 251 381 258 386
rect 251 379 253 381
rect 255 379 258 381
rect 240 370 245 377
rect 251 376 258 379
rect 260 388 268 390
rect 260 386 263 388
rect 265 386 268 388
rect 260 376 268 386
rect 270 383 275 390
rect 326 384 333 390
rect 270 380 278 383
rect 270 378 273 380
rect 275 378 278 380
rect 270 376 278 378
rect 273 373 278 376
rect 280 377 288 383
rect 280 375 283 377
rect 285 375 288 377
rect 280 373 288 375
rect 283 370 288 373
rect 290 381 297 383
rect 290 379 293 381
rect 295 379 297 381
rect 290 377 297 379
rect 315 381 322 384
rect 315 379 317 381
rect 319 379 322 381
rect 315 377 322 379
rect 290 370 295 377
rect 317 370 322 377
rect 324 374 333 384
rect 324 372 328 374
rect 330 372 333 374
rect 324 370 333 372
rect 335 370 340 390
rect 342 383 347 390
rect 353 388 360 390
rect 353 386 355 388
rect 357 386 360 388
rect 342 381 349 383
rect 342 379 345 381
rect 347 379 349 381
rect 342 377 349 379
rect 353 381 360 386
rect 353 379 355 381
rect 357 379 360 381
rect 342 370 347 377
rect 353 376 360 379
rect 362 388 370 390
rect 362 386 365 388
rect 367 386 370 388
rect 362 376 370 386
rect 372 383 377 390
rect 415 388 422 390
rect 415 386 417 388
rect 419 386 422 388
rect 372 380 380 383
rect 372 378 375 380
rect 377 378 380 380
rect 372 376 380 378
rect 375 373 380 376
rect 382 377 390 383
rect 382 375 385 377
rect 387 375 390 377
rect 382 373 390 375
rect 385 370 390 373
rect 392 381 399 383
rect 392 379 395 381
rect 397 379 399 381
rect 392 377 399 379
rect 415 381 422 386
rect 415 379 417 381
rect 419 379 422 381
rect 392 370 397 377
rect 415 376 422 379
rect 424 385 429 390
rect 437 385 442 387
rect 424 381 432 385
rect 424 379 427 381
rect 429 379 432 381
rect 424 377 432 379
rect 434 383 442 385
rect 434 381 437 383
rect 439 381 442 383
rect 434 379 442 381
rect 444 383 451 387
rect 479 384 486 390
rect 444 381 447 383
rect 449 381 451 383
rect 444 379 451 381
rect 468 381 475 384
rect 468 379 470 381
rect 472 379 475 381
rect 434 377 439 379
rect 424 376 429 377
rect 468 377 475 379
rect 470 370 475 377
rect 477 374 486 384
rect 477 372 481 374
rect 483 372 486 374
rect 477 370 486 372
rect 488 370 493 390
rect 495 383 500 390
rect 506 388 513 390
rect 506 386 508 388
rect 510 386 513 388
rect 495 381 502 383
rect 495 379 498 381
rect 500 379 502 381
rect 495 377 502 379
rect 506 381 513 386
rect 506 379 508 381
rect 510 379 513 381
rect 495 370 500 377
rect 506 376 513 379
rect 515 388 523 390
rect 515 386 518 388
rect 520 386 523 388
rect 515 376 523 386
rect 525 383 530 390
rect 580 384 587 390
rect 525 380 533 383
rect 525 378 528 380
rect 530 378 533 380
rect 525 376 533 378
rect 528 373 533 376
rect 535 377 543 383
rect 535 375 538 377
rect 540 375 543 377
rect 535 373 543 375
rect 538 370 543 373
rect 545 381 552 383
rect 545 379 548 381
rect 550 379 552 381
rect 545 377 552 379
rect 569 381 576 384
rect 569 379 571 381
rect 573 379 576 381
rect 569 377 576 379
rect 545 370 550 377
rect 571 370 576 377
rect 578 374 587 384
rect 578 372 582 374
rect 584 372 587 374
rect 578 370 587 372
rect 589 370 594 390
rect 596 383 601 390
rect 607 388 614 390
rect 607 386 609 388
rect 611 386 614 388
rect 596 381 603 383
rect 596 379 599 381
rect 601 379 603 381
rect 596 377 603 379
rect 607 381 614 386
rect 607 379 609 381
rect 611 379 614 381
rect 596 370 601 377
rect 607 376 614 379
rect 616 388 624 390
rect 616 386 619 388
rect 621 386 624 388
rect 616 376 624 386
rect 626 383 631 390
rect 679 384 686 390
rect 626 380 634 383
rect 626 378 629 380
rect 631 378 634 380
rect 626 376 634 378
rect 629 373 634 376
rect 636 377 644 383
rect 636 375 639 377
rect 641 375 644 377
rect 636 373 644 375
rect 639 370 644 373
rect 646 381 653 383
rect 646 379 649 381
rect 651 379 653 381
rect 646 377 653 379
rect 668 381 675 384
rect 668 379 670 381
rect 672 379 675 381
rect 668 377 675 379
rect 646 370 651 377
rect 670 370 675 377
rect 677 374 686 384
rect 677 372 681 374
rect 683 372 686 374
rect 677 370 686 372
rect 688 370 693 390
rect 695 383 700 390
rect 706 388 713 390
rect 706 386 708 388
rect 710 386 713 388
rect 695 381 702 383
rect 695 379 698 381
rect 700 379 702 381
rect 695 377 702 379
rect 706 381 713 386
rect 706 379 708 381
rect 710 379 713 381
rect 695 370 700 377
rect 706 376 713 379
rect 715 388 723 390
rect 715 386 718 388
rect 720 386 723 388
rect 715 376 723 386
rect 725 383 730 390
rect 725 380 733 383
rect 725 378 728 380
rect 730 378 733 380
rect 725 376 733 378
rect 728 373 733 376
rect 735 377 743 383
rect 735 375 738 377
rect 740 375 743 377
rect 735 373 743 375
rect 738 370 743 373
rect 745 381 752 383
rect 745 379 748 381
rect 750 379 752 381
rect 745 377 752 379
rect 745 370 750 377
rect 75 351 80 358
rect 73 349 80 351
rect 73 347 75 349
rect 77 347 80 349
rect 73 344 80 347
rect 82 356 91 358
rect 82 354 86 356
rect 88 354 91 356
rect 82 344 91 354
rect 84 338 91 344
rect 93 338 98 358
rect 100 351 105 358
rect 143 355 148 358
rect 133 352 138 355
rect 100 349 107 351
rect 100 347 103 349
rect 105 347 107 349
rect 100 345 107 347
rect 111 349 118 352
rect 111 347 113 349
rect 115 347 118 349
rect 100 338 105 345
rect 111 342 118 347
rect 111 340 113 342
rect 115 340 118 342
rect 111 338 118 340
rect 120 342 128 352
rect 120 340 123 342
rect 125 340 128 342
rect 120 338 128 340
rect 130 350 138 352
rect 130 348 133 350
rect 135 348 138 350
rect 130 345 138 348
rect 140 353 148 355
rect 140 351 143 353
rect 145 351 148 353
rect 140 345 148 351
rect 150 351 155 358
rect 150 349 157 351
rect 150 347 153 349
rect 155 347 157 349
rect 150 345 157 347
rect 161 349 168 352
rect 161 347 163 349
rect 165 347 168 349
rect 130 338 135 345
rect 161 342 168 347
rect 161 340 163 342
rect 165 340 168 342
rect 161 338 168 340
rect 170 351 175 352
rect 170 349 178 351
rect 170 347 173 349
rect 175 347 178 349
rect 170 343 178 347
rect 180 349 185 351
rect 216 351 221 358
rect 214 349 221 351
rect 180 347 188 349
rect 180 345 183 347
rect 185 345 188 347
rect 180 343 188 345
rect 170 338 175 343
rect 183 341 188 343
rect 190 347 197 349
rect 190 345 193 347
rect 195 345 197 347
rect 190 341 197 345
rect 214 347 216 349
rect 218 347 221 349
rect 214 344 221 347
rect 223 356 232 358
rect 223 354 227 356
rect 229 354 232 356
rect 223 344 232 354
rect 225 338 232 344
rect 234 338 239 358
rect 241 351 246 358
rect 284 355 289 358
rect 274 352 279 355
rect 241 349 248 351
rect 241 347 244 349
rect 246 347 248 349
rect 241 345 248 347
rect 252 349 259 352
rect 252 347 254 349
rect 256 347 259 349
rect 241 338 246 345
rect 252 342 259 347
rect 252 340 254 342
rect 256 340 259 342
rect 252 338 259 340
rect 261 342 269 352
rect 261 340 264 342
rect 266 340 269 342
rect 261 338 269 340
rect 271 350 279 352
rect 271 348 274 350
rect 276 348 279 350
rect 271 345 279 348
rect 281 353 289 355
rect 281 351 284 353
rect 286 351 289 353
rect 281 345 289 351
rect 291 351 296 358
rect 316 351 321 358
rect 291 349 298 351
rect 291 347 294 349
rect 296 347 298 349
rect 291 345 298 347
rect 314 349 321 351
rect 314 347 316 349
rect 318 347 321 349
rect 314 345 321 347
rect 323 355 328 358
rect 323 353 331 355
rect 323 351 326 353
rect 328 351 331 353
rect 323 345 331 351
rect 333 352 338 355
rect 333 350 341 352
rect 333 348 336 350
rect 338 348 341 350
rect 333 345 341 348
rect 271 338 276 345
rect 336 338 341 345
rect 343 342 351 352
rect 343 340 346 342
rect 348 340 351 342
rect 343 338 351 340
rect 353 349 360 352
rect 366 351 371 358
rect 353 347 356 349
rect 358 347 360 349
rect 353 342 360 347
rect 364 349 371 351
rect 364 347 366 349
rect 368 347 371 349
rect 364 345 371 347
rect 353 340 356 342
rect 358 340 360 342
rect 353 338 360 340
rect 366 338 371 345
rect 373 338 378 358
rect 380 356 389 358
rect 380 354 383 356
rect 385 354 389 356
rect 380 344 389 354
rect 391 351 396 358
rect 391 349 398 351
rect 391 347 394 349
rect 396 347 398 349
rect 391 344 398 347
rect 415 349 422 352
rect 415 347 417 349
rect 419 347 422 349
rect 380 338 387 344
rect 415 342 422 347
rect 415 340 417 342
rect 419 340 422 342
rect 415 338 422 340
rect 424 351 429 352
rect 424 349 432 351
rect 424 347 427 349
rect 429 347 432 349
rect 424 343 432 347
rect 434 349 439 351
rect 470 351 475 358
rect 468 349 475 351
rect 434 347 442 349
rect 434 345 437 347
rect 439 345 442 347
rect 434 343 442 345
rect 424 338 429 343
rect 437 341 442 343
rect 444 347 451 349
rect 444 345 447 347
rect 449 345 451 347
rect 444 341 451 345
rect 468 347 470 349
rect 472 347 475 349
rect 468 344 475 347
rect 477 356 486 358
rect 477 354 481 356
rect 483 354 486 356
rect 477 344 486 354
rect 479 338 486 344
rect 488 338 493 358
rect 495 351 500 358
rect 538 355 543 358
rect 528 352 533 355
rect 495 349 502 351
rect 495 347 498 349
rect 500 347 502 349
rect 495 345 502 347
rect 506 349 513 352
rect 506 347 508 349
rect 510 347 513 349
rect 495 338 500 345
rect 506 342 513 347
rect 506 340 508 342
rect 510 340 513 342
rect 506 338 513 340
rect 515 342 523 352
rect 515 340 518 342
rect 520 340 523 342
rect 515 338 523 340
rect 525 350 533 352
rect 525 348 528 350
rect 530 348 533 350
rect 525 345 533 348
rect 535 353 543 355
rect 535 351 538 353
rect 540 351 543 353
rect 535 345 543 351
rect 545 351 550 358
rect 571 351 576 358
rect 545 349 552 351
rect 545 347 548 349
rect 550 347 552 349
rect 545 345 552 347
rect 569 349 576 351
rect 569 347 571 349
rect 573 347 576 349
rect 525 338 530 345
rect 569 344 576 347
rect 578 356 587 358
rect 578 354 582 356
rect 584 354 587 356
rect 578 344 587 354
rect 580 338 587 344
rect 589 338 594 358
rect 596 351 601 358
rect 639 355 644 358
rect 629 352 634 355
rect 596 349 603 351
rect 596 347 599 349
rect 601 347 603 349
rect 596 345 603 347
rect 607 349 614 352
rect 607 347 609 349
rect 611 347 614 349
rect 596 338 601 345
rect 607 342 614 347
rect 607 340 609 342
rect 611 340 614 342
rect 607 338 614 340
rect 616 342 624 352
rect 616 340 619 342
rect 621 340 624 342
rect 616 338 624 340
rect 626 350 634 352
rect 626 348 629 350
rect 631 348 634 350
rect 626 345 634 348
rect 636 353 644 355
rect 636 351 639 353
rect 641 351 644 353
rect 636 345 644 351
rect 646 351 651 358
rect 670 351 675 358
rect 646 349 653 351
rect 646 347 649 349
rect 651 347 653 349
rect 646 345 653 347
rect 668 349 675 351
rect 668 347 670 349
rect 672 347 675 349
rect 626 338 631 345
rect 668 344 675 347
rect 677 356 686 358
rect 677 354 681 356
rect 683 354 686 356
rect 677 344 686 354
rect 679 338 686 344
rect 688 338 693 358
rect 695 351 700 358
rect 738 355 743 358
rect 728 352 733 355
rect 695 349 702 351
rect 695 347 698 349
rect 700 347 702 349
rect 695 345 702 347
rect 706 349 713 352
rect 706 347 708 349
rect 710 347 713 349
rect 695 338 700 345
rect 706 342 713 347
rect 706 340 708 342
rect 710 340 713 342
rect 706 338 713 340
rect 715 342 723 352
rect 715 340 718 342
rect 720 340 723 342
rect 715 338 723 340
rect 725 350 733 352
rect 725 348 728 350
rect 730 348 733 350
rect 725 345 733 348
rect 735 353 743 355
rect 735 351 738 353
rect 740 351 743 353
rect 735 345 743 351
rect 745 351 750 358
rect 745 349 752 351
rect 745 347 748 349
rect 750 347 752 349
rect 745 345 752 347
rect 725 338 730 345
rect 71 244 78 246
rect 71 242 73 244
rect 75 242 78 244
rect 71 237 78 242
rect 71 235 73 237
rect 75 235 78 237
rect 71 232 78 235
rect 80 241 85 246
rect 93 241 98 243
rect 80 237 88 241
rect 80 235 83 237
rect 85 235 88 237
rect 80 233 88 235
rect 90 239 98 241
rect 90 237 93 239
rect 95 237 98 239
rect 90 235 98 237
rect 100 239 107 243
rect 123 240 130 246
rect 100 237 103 239
rect 105 237 107 239
rect 100 235 107 237
rect 112 237 119 240
rect 112 235 114 237
rect 116 235 119 237
rect 90 233 95 235
rect 80 232 85 233
rect 112 233 119 235
rect 114 226 119 233
rect 121 230 130 240
rect 121 228 125 230
rect 127 228 130 230
rect 121 226 130 228
rect 132 226 137 246
rect 139 239 144 246
rect 150 244 157 246
rect 150 242 152 244
rect 154 242 157 244
rect 139 237 146 239
rect 139 235 142 237
rect 144 235 146 237
rect 139 233 146 235
rect 150 237 157 242
rect 150 235 152 237
rect 154 235 157 237
rect 139 226 144 233
rect 150 232 157 235
rect 159 244 167 246
rect 159 242 162 244
rect 164 242 167 244
rect 159 232 167 242
rect 169 239 174 246
rect 224 240 231 246
rect 169 236 177 239
rect 169 234 172 236
rect 174 234 177 236
rect 169 232 177 234
rect 172 229 177 232
rect 179 233 187 239
rect 179 231 182 233
rect 184 231 187 233
rect 179 229 187 231
rect 182 226 187 229
rect 189 237 196 239
rect 189 235 192 237
rect 194 235 196 237
rect 189 233 196 235
rect 213 237 220 240
rect 213 235 215 237
rect 217 235 220 237
rect 213 233 220 235
rect 189 226 194 233
rect 215 226 220 233
rect 222 230 231 240
rect 222 228 226 230
rect 228 228 231 230
rect 222 226 231 228
rect 233 226 238 246
rect 240 239 245 246
rect 251 244 258 246
rect 251 242 253 244
rect 255 242 258 244
rect 240 237 247 239
rect 240 235 243 237
rect 245 235 247 237
rect 240 233 247 235
rect 251 237 258 242
rect 251 235 253 237
rect 255 235 258 237
rect 240 226 245 233
rect 251 232 258 235
rect 260 244 268 246
rect 260 242 263 244
rect 265 242 268 244
rect 260 232 268 242
rect 270 239 275 246
rect 325 240 332 246
rect 270 236 278 239
rect 270 234 273 236
rect 275 234 278 236
rect 270 232 278 234
rect 273 229 278 232
rect 280 233 288 239
rect 280 231 283 233
rect 285 231 288 233
rect 280 229 288 231
rect 283 226 288 229
rect 290 237 297 239
rect 290 235 293 237
rect 295 235 297 237
rect 290 233 297 235
rect 314 237 321 240
rect 314 235 316 237
rect 318 235 321 237
rect 314 233 321 235
rect 290 226 295 233
rect 316 226 321 233
rect 323 230 332 240
rect 323 228 327 230
rect 329 228 332 230
rect 323 226 332 228
rect 334 226 339 246
rect 341 239 346 246
rect 352 244 359 246
rect 352 242 354 244
rect 356 242 359 244
rect 341 237 348 239
rect 341 235 344 237
rect 346 235 348 237
rect 341 233 348 235
rect 352 237 359 242
rect 352 235 354 237
rect 356 235 359 237
rect 341 226 346 233
rect 352 232 359 235
rect 361 244 369 246
rect 361 242 364 244
rect 366 242 369 244
rect 361 232 369 242
rect 371 239 376 246
rect 414 244 421 246
rect 414 242 416 244
rect 418 242 421 244
rect 371 236 379 239
rect 371 234 374 236
rect 376 234 379 236
rect 371 232 379 234
rect 374 229 379 232
rect 381 233 389 239
rect 381 231 384 233
rect 386 231 389 233
rect 381 229 389 231
rect 384 226 389 229
rect 391 237 398 239
rect 391 235 394 237
rect 396 235 398 237
rect 391 233 398 235
rect 414 237 421 242
rect 414 235 416 237
rect 418 235 421 237
rect 391 226 396 233
rect 414 232 421 235
rect 423 241 428 246
rect 436 241 441 243
rect 423 237 431 241
rect 423 235 426 237
rect 428 235 431 237
rect 423 233 431 235
rect 433 239 441 241
rect 433 237 436 239
rect 438 237 441 239
rect 433 235 441 237
rect 443 239 450 243
rect 478 240 485 246
rect 443 237 446 239
rect 448 237 450 239
rect 443 235 450 237
rect 467 237 474 240
rect 467 235 469 237
rect 471 235 474 237
rect 433 233 438 235
rect 423 232 428 233
rect 467 233 474 235
rect 469 226 474 233
rect 476 230 485 240
rect 476 228 480 230
rect 482 228 485 230
rect 476 226 485 228
rect 487 226 492 246
rect 494 239 499 246
rect 505 244 512 246
rect 505 242 507 244
rect 509 242 512 244
rect 494 237 501 239
rect 494 235 497 237
rect 499 235 501 237
rect 494 233 501 235
rect 505 237 512 242
rect 505 235 507 237
rect 509 235 512 237
rect 494 226 499 233
rect 505 232 512 235
rect 514 244 522 246
rect 514 242 517 244
rect 519 242 522 244
rect 514 232 522 242
rect 524 239 529 246
rect 579 240 586 246
rect 524 236 532 239
rect 524 234 527 236
rect 529 234 532 236
rect 524 232 532 234
rect 527 229 532 232
rect 534 233 542 239
rect 534 231 537 233
rect 539 231 542 233
rect 534 229 542 231
rect 537 226 542 229
rect 544 237 551 239
rect 544 235 547 237
rect 549 235 551 237
rect 544 233 551 235
rect 568 237 575 240
rect 568 235 570 237
rect 572 235 575 237
rect 568 233 575 235
rect 544 226 549 233
rect 570 226 575 233
rect 577 230 586 240
rect 577 228 581 230
rect 583 228 586 230
rect 577 226 586 228
rect 588 226 593 246
rect 595 239 600 246
rect 606 244 613 246
rect 606 242 608 244
rect 610 242 613 244
rect 595 237 602 239
rect 595 235 598 237
rect 600 235 602 237
rect 595 233 602 235
rect 606 237 613 242
rect 606 235 608 237
rect 610 235 613 237
rect 595 226 600 233
rect 606 232 613 235
rect 615 244 623 246
rect 615 242 618 244
rect 620 242 623 244
rect 615 232 623 242
rect 625 239 630 246
rect 678 240 685 246
rect 625 236 633 239
rect 625 234 628 236
rect 630 234 633 236
rect 625 232 633 234
rect 628 229 633 232
rect 635 233 643 239
rect 635 231 638 233
rect 640 231 643 233
rect 635 229 643 231
rect 638 226 643 229
rect 645 237 652 239
rect 645 235 648 237
rect 650 235 652 237
rect 645 233 652 235
rect 667 237 674 240
rect 667 235 669 237
rect 671 235 674 237
rect 667 233 674 235
rect 645 226 650 233
rect 669 226 674 233
rect 676 230 685 240
rect 676 228 680 230
rect 682 228 685 230
rect 676 226 685 228
rect 687 226 692 246
rect 694 239 699 246
rect 705 244 712 246
rect 705 242 707 244
rect 709 242 712 244
rect 694 237 701 239
rect 694 235 697 237
rect 699 235 701 237
rect 694 233 701 235
rect 705 237 712 242
rect 705 235 707 237
rect 709 235 712 237
rect 694 226 699 233
rect 705 232 712 235
rect 714 244 722 246
rect 714 242 717 244
rect 719 242 722 244
rect 714 232 722 242
rect 724 239 729 246
rect 724 236 732 239
rect 724 234 727 236
rect 729 234 732 236
rect 724 232 732 234
rect 727 229 732 232
rect 734 233 742 239
rect 734 231 737 233
rect 739 231 742 233
rect 734 229 742 231
rect 737 226 742 229
rect 744 237 751 239
rect 744 235 747 237
rect 749 235 751 237
rect 744 233 751 235
rect 744 226 749 233
<< pdif >>
rect 71 572 78 574
rect 71 570 73 572
rect 75 570 78 572
rect 71 565 78 570
rect 71 563 73 565
rect 75 563 78 565
rect 71 555 78 563
rect 80 566 88 574
rect 80 564 83 566
rect 85 564 88 566
rect 80 559 88 564
rect 80 557 83 559
rect 85 557 88 559
rect 80 555 88 557
rect 90 572 98 574
rect 90 570 93 572
rect 95 570 98 572
rect 90 565 98 570
rect 90 563 93 565
rect 95 563 98 565
rect 90 555 98 563
rect 92 546 98 555
rect 100 567 105 574
rect 111 572 118 574
rect 111 570 113 572
rect 115 570 118 572
rect 100 565 107 567
rect 100 563 103 565
rect 105 563 107 565
rect 100 558 107 563
rect 100 556 103 558
rect 105 556 107 558
rect 100 554 107 556
rect 111 565 118 570
rect 111 563 113 565
rect 115 563 118 565
rect 111 555 118 563
rect 120 566 128 574
rect 120 564 123 566
rect 125 564 128 566
rect 120 559 128 564
rect 120 557 123 559
rect 125 557 128 559
rect 120 555 128 557
rect 130 572 138 574
rect 130 570 133 572
rect 135 570 138 572
rect 130 565 138 570
rect 130 563 133 565
rect 135 563 138 565
rect 130 555 138 563
rect 100 546 105 554
rect 132 546 138 555
rect 140 567 145 574
rect 140 565 147 567
rect 140 563 143 565
rect 145 563 147 565
rect 140 558 147 563
rect 154 559 159 574
rect 140 556 143 558
rect 145 556 147 558
rect 140 554 147 556
rect 152 557 159 559
rect 152 555 154 557
rect 156 555 159 557
rect 140 546 145 554
rect 152 550 159 555
rect 152 548 154 550
rect 156 548 159 550
rect 152 546 159 548
rect 161 572 169 574
rect 161 570 164 572
rect 166 570 169 572
rect 161 565 169 570
rect 161 563 164 565
rect 166 563 169 565
rect 161 546 169 563
rect 171 564 179 574
rect 171 562 174 564
rect 176 562 179 564
rect 171 557 179 562
rect 171 555 174 557
rect 176 555 179 557
rect 171 546 179 555
rect 181 572 195 574
rect 181 570 186 572
rect 188 571 195 572
rect 218 572 227 574
rect 188 570 197 571
rect 181 565 197 570
rect 181 563 186 565
rect 188 563 197 565
rect 181 546 197 563
rect 199 546 204 571
rect 206 562 211 571
rect 218 570 221 572
rect 223 570 227 572
rect 218 562 227 570
rect 206 553 214 562
rect 206 551 209 553
rect 211 551 214 553
rect 206 549 214 551
rect 216 549 227 562
rect 229 562 234 574
rect 250 562 255 574
rect 229 560 236 562
rect 229 558 232 560
rect 234 558 236 560
rect 229 553 236 558
rect 229 551 232 553
rect 234 551 236 553
rect 229 549 236 551
rect 248 560 255 562
rect 248 558 250 560
rect 252 558 255 560
rect 248 553 255 558
rect 248 551 250 553
rect 252 551 255 553
rect 248 549 255 551
rect 257 572 266 574
rect 257 570 261 572
rect 263 570 266 572
rect 289 572 303 574
rect 289 571 296 572
rect 257 562 266 570
rect 273 562 278 571
rect 257 549 268 562
rect 270 553 278 562
rect 270 551 273 553
rect 275 551 278 553
rect 270 549 278 551
rect 206 546 211 549
rect 273 546 278 549
rect 280 546 285 571
rect 287 570 296 571
rect 298 570 303 572
rect 287 565 303 570
rect 287 563 296 565
rect 298 563 303 565
rect 287 546 303 563
rect 305 564 313 574
rect 305 562 308 564
rect 310 562 313 564
rect 305 557 313 562
rect 305 555 308 557
rect 310 555 313 557
rect 305 546 313 555
rect 315 572 323 574
rect 315 570 318 572
rect 320 570 323 572
rect 315 565 323 570
rect 315 563 318 565
rect 320 563 323 565
rect 315 546 323 563
rect 325 559 330 574
rect 339 567 344 574
rect 337 565 344 567
rect 337 563 339 565
rect 341 563 344 565
rect 325 557 332 559
rect 325 555 328 557
rect 330 555 332 557
rect 325 550 332 555
rect 337 558 344 563
rect 337 556 339 558
rect 341 556 344 558
rect 337 554 344 556
rect 325 548 328 550
rect 330 548 332 550
rect 325 546 332 548
rect 339 546 344 554
rect 346 572 354 574
rect 346 570 349 572
rect 351 570 354 572
rect 346 565 354 570
rect 346 563 349 565
rect 351 563 354 565
rect 346 555 354 563
rect 356 566 364 574
rect 356 564 359 566
rect 361 564 364 566
rect 356 559 364 564
rect 356 557 359 559
rect 361 557 364 559
rect 356 555 364 557
rect 366 572 373 574
rect 366 570 369 572
rect 371 570 373 572
rect 366 565 373 570
rect 379 567 384 574
rect 366 563 369 565
rect 371 563 373 565
rect 366 555 373 563
rect 377 565 384 567
rect 377 563 379 565
rect 381 563 384 565
rect 377 558 384 563
rect 377 556 379 558
rect 381 556 384 558
rect 346 546 352 555
rect 377 554 384 556
rect 379 546 384 554
rect 386 572 394 574
rect 386 570 389 572
rect 391 570 394 572
rect 386 565 394 570
rect 386 563 389 565
rect 391 563 394 565
rect 386 555 394 563
rect 396 566 404 574
rect 396 564 399 566
rect 401 564 404 566
rect 396 559 404 564
rect 396 557 399 559
rect 401 557 404 559
rect 396 555 404 557
rect 406 572 413 574
rect 406 570 409 572
rect 411 570 413 572
rect 406 565 413 570
rect 406 563 409 565
rect 411 563 413 565
rect 406 555 413 563
rect 420 562 425 574
rect 418 560 425 562
rect 418 558 420 560
rect 422 558 425 560
rect 386 546 392 555
rect 418 553 425 558
rect 418 551 420 553
rect 422 551 425 553
rect 418 549 425 551
rect 427 572 436 574
rect 427 570 431 572
rect 433 570 436 572
rect 459 572 473 574
rect 459 571 466 572
rect 427 562 436 570
rect 443 562 448 571
rect 427 549 438 562
rect 440 553 448 562
rect 440 551 443 553
rect 445 551 448 553
rect 440 549 448 551
rect 443 546 448 549
rect 450 546 455 571
rect 457 570 466 571
rect 468 570 473 572
rect 457 565 473 570
rect 457 563 466 565
rect 468 563 473 565
rect 457 546 473 563
rect 475 564 483 574
rect 475 562 478 564
rect 480 562 483 564
rect 475 557 483 562
rect 475 555 478 557
rect 480 555 483 557
rect 475 546 483 555
rect 485 572 493 574
rect 485 570 488 572
rect 490 570 493 572
rect 485 565 493 570
rect 485 563 488 565
rect 490 563 493 565
rect 485 546 493 563
rect 495 559 500 574
rect 509 567 514 574
rect 507 565 514 567
rect 507 563 509 565
rect 511 563 514 565
rect 495 557 502 559
rect 495 555 498 557
rect 500 555 502 557
rect 495 550 502 555
rect 507 558 514 563
rect 507 556 509 558
rect 511 556 514 558
rect 507 554 514 556
rect 495 548 498 550
rect 500 548 502 550
rect 495 546 502 548
rect 509 546 514 554
rect 516 572 524 574
rect 516 570 519 572
rect 521 570 524 572
rect 516 565 524 570
rect 516 563 519 565
rect 521 563 524 565
rect 516 555 524 563
rect 526 566 534 574
rect 526 564 529 566
rect 531 564 534 566
rect 526 559 534 564
rect 526 557 529 559
rect 531 557 534 559
rect 526 555 534 557
rect 536 572 543 574
rect 536 570 539 572
rect 541 570 543 572
rect 536 565 543 570
rect 549 567 554 574
rect 536 563 539 565
rect 541 563 543 565
rect 536 555 543 563
rect 547 565 554 567
rect 547 563 549 565
rect 551 563 554 565
rect 547 558 554 563
rect 547 556 549 558
rect 551 556 554 558
rect 516 546 522 555
rect 547 554 554 556
rect 549 546 554 554
rect 556 572 564 574
rect 556 570 559 572
rect 561 570 564 572
rect 556 565 564 570
rect 556 563 559 565
rect 561 563 564 565
rect 556 555 564 563
rect 566 566 574 574
rect 566 564 569 566
rect 571 564 574 566
rect 566 559 574 564
rect 566 557 569 559
rect 571 557 574 559
rect 566 555 574 557
rect 576 572 583 574
rect 576 570 579 572
rect 581 570 583 572
rect 576 565 583 570
rect 576 563 579 565
rect 581 563 583 565
rect 576 555 583 563
rect 587 572 594 574
rect 587 570 589 572
rect 591 570 594 572
rect 587 565 594 570
rect 587 563 589 565
rect 591 563 594 565
rect 587 555 594 563
rect 596 566 604 574
rect 596 564 599 566
rect 601 564 604 566
rect 596 559 604 564
rect 596 557 599 559
rect 601 557 604 559
rect 596 555 604 557
rect 606 572 614 574
rect 606 570 609 572
rect 611 570 614 572
rect 606 565 614 570
rect 606 563 609 565
rect 611 563 614 565
rect 606 555 614 563
rect 556 546 562 555
rect 608 546 614 555
rect 616 567 621 574
rect 627 572 634 574
rect 627 570 629 572
rect 631 570 634 572
rect 616 565 623 567
rect 616 563 619 565
rect 621 563 623 565
rect 616 558 623 563
rect 616 556 619 558
rect 621 556 623 558
rect 616 554 623 556
rect 627 565 634 570
rect 627 563 629 565
rect 631 563 634 565
rect 627 555 634 563
rect 636 566 644 574
rect 636 564 639 566
rect 641 564 644 566
rect 636 559 644 564
rect 636 557 639 559
rect 641 557 644 559
rect 636 555 644 557
rect 646 572 654 574
rect 646 570 649 572
rect 651 570 654 572
rect 646 565 654 570
rect 646 563 649 565
rect 651 563 654 565
rect 646 555 654 563
rect 616 546 621 554
rect 648 546 654 555
rect 656 567 661 574
rect 656 565 663 567
rect 656 563 659 565
rect 661 563 663 565
rect 656 558 663 563
rect 670 559 675 574
rect 656 556 659 558
rect 661 556 663 558
rect 656 554 663 556
rect 668 557 675 559
rect 668 555 670 557
rect 672 555 675 557
rect 656 546 661 554
rect 668 550 675 555
rect 668 548 670 550
rect 672 548 675 550
rect 668 546 675 548
rect 677 572 685 574
rect 677 570 680 572
rect 682 570 685 572
rect 677 565 685 570
rect 677 563 680 565
rect 682 563 685 565
rect 677 546 685 563
rect 687 564 695 574
rect 687 562 690 564
rect 692 562 695 564
rect 687 557 695 562
rect 687 555 690 557
rect 692 555 695 557
rect 687 546 695 555
rect 697 572 711 574
rect 697 570 702 572
rect 704 571 711 572
rect 734 572 743 574
rect 704 570 713 571
rect 697 565 713 570
rect 697 563 702 565
rect 704 563 713 565
rect 697 546 713 563
rect 715 546 720 571
rect 722 562 727 571
rect 734 570 737 572
rect 739 570 743 572
rect 734 562 743 570
rect 722 553 730 562
rect 722 551 725 553
rect 727 551 730 553
rect 722 549 730 551
rect 732 549 743 562
rect 745 562 750 574
rect 745 560 752 562
rect 745 558 748 560
rect 750 558 752 560
rect 745 553 752 558
rect 745 551 748 553
rect 750 551 752 553
rect 745 549 752 551
rect 722 546 727 549
rect 92 461 98 470
rect 71 453 78 461
rect 71 451 73 453
rect 75 451 78 453
rect 71 446 78 451
rect 71 444 73 446
rect 75 444 78 446
rect 71 442 78 444
rect 80 459 88 461
rect 80 457 83 459
rect 85 457 88 459
rect 80 452 88 457
rect 80 450 83 452
rect 85 450 88 452
rect 80 442 88 450
rect 90 453 98 461
rect 90 451 93 453
rect 95 451 98 453
rect 90 446 98 451
rect 90 444 93 446
rect 95 444 98 446
rect 90 442 98 444
rect 100 462 105 470
rect 100 460 107 462
rect 132 461 138 470
rect 100 458 103 460
rect 105 458 107 460
rect 100 453 107 458
rect 100 451 103 453
rect 105 451 107 453
rect 100 449 107 451
rect 111 453 118 461
rect 111 451 113 453
rect 115 451 118 453
rect 100 442 105 449
rect 111 446 118 451
rect 111 444 113 446
rect 115 444 118 446
rect 111 442 118 444
rect 120 459 128 461
rect 120 457 123 459
rect 125 457 128 459
rect 120 452 128 457
rect 120 450 123 452
rect 125 450 128 452
rect 120 442 128 450
rect 130 453 138 461
rect 130 451 133 453
rect 135 451 138 453
rect 130 446 138 451
rect 130 444 133 446
rect 135 444 138 446
rect 130 442 138 444
rect 140 462 145 470
rect 152 468 159 470
rect 152 466 154 468
rect 156 466 159 468
rect 140 460 147 462
rect 140 458 143 460
rect 145 458 147 460
rect 140 453 147 458
rect 152 457 159 466
rect 140 451 143 453
rect 145 451 147 453
rect 140 449 147 451
rect 140 442 145 449
rect 154 442 159 457
rect 161 453 169 470
rect 161 451 164 453
rect 166 451 169 453
rect 161 446 169 451
rect 161 444 164 446
rect 166 444 169 446
rect 161 442 169 444
rect 171 461 179 470
rect 171 459 174 461
rect 176 459 179 461
rect 171 454 179 459
rect 171 452 174 454
rect 176 452 179 454
rect 171 442 179 452
rect 181 453 197 470
rect 181 451 186 453
rect 188 451 197 453
rect 181 446 197 451
rect 181 444 186 446
rect 188 445 197 446
rect 199 445 204 470
rect 206 467 211 470
rect 273 467 278 470
rect 206 465 214 467
rect 206 463 209 465
rect 211 463 214 465
rect 206 454 214 463
rect 216 454 227 467
rect 206 445 211 454
rect 218 446 227 454
rect 188 444 195 445
rect 181 442 195 444
rect 218 444 221 446
rect 223 444 227 446
rect 218 442 227 444
rect 229 465 236 467
rect 229 463 232 465
rect 234 463 236 465
rect 229 458 236 463
rect 229 456 232 458
rect 234 456 236 458
rect 229 454 236 456
rect 248 465 255 467
rect 248 463 250 465
rect 252 463 255 465
rect 248 458 255 463
rect 248 456 250 458
rect 252 456 255 458
rect 248 454 255 456
rect 229 442 234 454
rect 250 442 255 454
rect 257 454 268 467
rect 270 465 278 467
rect 270 463 273 465
rect 275 463 278 465
rect 270 454 278 463
rect 257 446 266 454
rect 257 444 261 446
rect 263 444 266 446
rect 273 445 278 454
rect 280 445 285 470
rect 287 453 303 470
rect 287 451 296 453
rect 298 451 303 453
rect 287 446 303 451
rect 287 445 296 446
rect 257 442 266 444
rect 289 444 296 445
rect 298 444 303 446
rect 289 442 303 444
rect 305 461 313 470
rect 305 459 308 461
rect 310 459 313 461
rect 305 454 313 459
rect 305 452 308 454
rect 310 452 313 454
rect 305 442 313 452
rect 315 453 323 470
rect 315 451 318 453
rect 320 451 323 453
rect 315 446 323 451
rect 315 444 318 446
rect 320 444 323 446
rect 315 442 323 444
rect 325 468 332 470
rect 325 466 328 468
rect 330 466 332 468
rect 325 461 332 466
rect 339 462 344 470
rect 325 459 328 461
rect 330 459 332 461
rect 325 457 332 459
rect 337 460 344 462
rect 337 458 339 460
rect 341 458 344 460
rect 325 442 330 457
rect 337 453 344 458
rect 337 451 339 453
rect 341 451 344 453
rect 337 449 344 451
rect 339 442 344 449
rect 346 461 352 470
rect 379 462 384 470
rect 346 453 354 461
rect 346 451 349 453
rect 351 451 354 453
rect 346 446 354 451
rect 346 444 349 446
rect 351 444 354 446
rect 346 442 354 444
rect 356 459 364 461
rect 356 457 359 459
rect 361 457 364 459
rect 356 452 364 457
rect 356 450 359 452
rect 361 450 364 452
rect 356 442 364 450
rect 366 453 373 461
rect 366 451 369 453
rect 371 451 373 453
rect 366 446 373 451
rect 377 460 384 462
rect 377 458 379 460
rect 381 458 384 460
rect 377 453 384 458
rect 377 451 379 453
rect 381 451 384 453
rect 377 449 384 451
rect 366 444 369 446
rect 371 444 373 446
rect 366 442 373 444
rect 379 442 384 449
rect 386 461 392 470
rect 443 467 448 470
rect 418 465 425 467
rect 418 463 420 465
rect 422 463 425 465
rect 386 453 394 461
rect 386 451 389 453
rect 391 451 394 453
rect 386 446 394 451
rect 386 444 389 446
rect 391 444 394 446
rect 386 442 394 444
rect 396 459 404 461
rect 396 457 399 459
rect 401 457 404 459
rect 396 452 404 457
rect 396 450 399 452
rect 401 450 404 452
rect 396 442 404 450
rect 406 453 413 461
rect 418 458 425 463
rect 418 456 420 458
rect 422 456 425 458
rect 418 454 425 456
rect 406 451 409 453
rect 411 451 413 453
rect 406 446 413 451
rect 406 444 409 446
rect 411 444 413 446
rect 406 442 413 444
rect 420 442 425 454
rect 427 454 438 467
rect 440 465 448 467
rect 440 463 443 465
rect 445 463 448 465
rect 440 454 448 463
rect 427 446 436 454
rect 427 444 431 446
rect 433 444 436 446
rect 443 445 448 454
rect 450 445 455 470
rect 457 453 473 470
rect 457 451 466 453
rect 468 451 473 453
rect 457 446 473 451
rect 457 445 466 446
rect 427 442 436 444
rect 459 444 466 445
rect 468 444 473 446
rect 459 442 473 444
rect 475 461 483 470
rect 475 459 478 461
rect 480 459 483 461
rect 475 454 483 459
rect 475 452 478 454
rect 480 452 483 454
rect 475 442 483 452
rect 485 453 493 470
rect 485 451 488 453
rect 490 451 493 453
rect 485 446 493 451
rect 485 444 488 446
rect 490 444 493 446
rect 485 442 493 444
rect 495 468 502 470
rect 495 466 498 468
rect 500 466 502 468
rect 495 461 502 466
rect 509 462 514 470
rect 495 459 498 461
rect 500 459 502 461
rect 495 457 502 459
rect 507 460 514 462
rect 507 458 509 460
rect 511 458 514 460
rect 495 442 500 457
rect 507 453 514 458
rect 507 451 509 453
rect 511 451 514 453
rect 507 449 514 451
rect 509 442 514 449
rect 516 461 522 470
rect 549 462 554 470
rect 516 453 524 461
rect 516 451 519 453
rect 521 451 524 453
rect 516 446 524 451
rect 516 444 519 446
rect 521 444 524 446
rect 516 442 524 444
rect 526 459 534 461
rect 526 457 529 459
rect 531 457 534 459
rect 526 452 534 457
rect 526 450 529 452
rect 531 450 534 452
rect 526 442 534 450
rect 536 453 543 461
rect 536 451 539 453
rect 541 451 543 453
rect 536 446 543 451
rect 547 460 554 462
rect 547 458 549 460
rect 551 458 554 460
rect 547 453 554 458
rect 547 451 549 453
rect 551 451 554 453
rect 547 449 554 451
rect 536 444 539 446
rect 541 444 543 446
rect 536 442 543 444
rect 549 442 554 449
rect 556 461 562 470
rect 608 461 614 470
rect 556 453 564 461
rect 556 451 559 453
rect 561 451 564 453
rect 556 446 564 451
rect 556 444 559 446
rect 561 444 564 446
rect 556 442 564 444
rect 566 459 574 461
rect 566 457 569 459
rect 571 457 574 459
rect 566 452 574 457
rect 566 450 569 452
rect 571 450 574 452
rect 566 442 574 450
rect 576 453 583 461
rect 576 451 579 453
rect 581 451 583 453
rect 576 446 583 451
rect 576 444 579 446
rect 581 444 583 446
rect 576 442 583 444
rect 587 453 594 461
rect 587 451 589 453
rect 591 451 594 453
rect 587 446 594 451
rect 587 444 589 446
rect 591 444 594 446
rect 587 442 594 444
rect 596 459 604 461
rect 596 457 599 459
rect 601 457 604 459
rect 596 452 604 457
rect 596 450 599 452
rect 601 450 604 452
rect 596 442 604 450
rect 606 453 614 461
rect 606 451 609 453
rect 611 451 614 453
rect 606 446 614 451
rect 606 444 609 446
rect 611 444 614 446
rect 606 442 614 444
rect 616 462 621 470
rect 616 460 623 462
rect 648 461 654 470
rect 616 458 619 460
rect 621 458 623 460
rect 616 453 623 458
rect 616 451 619 453
rect 621 451 623 453
rect 616 449 623 451
rect 627 453 634 461
rect 627 451 629 453
rect 631 451 634 453
rect 616 442 621 449
rect 627 446 634 451
rect 627 444 629 446
rect 631 444 634 446
rect 627 442 634 444
rect 636 459 644 461
rect 636 457 639 459
rect 641 457 644 459
rect 636 452 644 457
rect 636 450 639 452
rect 641 450 644 452
rect 636 442 644 450
rect 646 453 654 461
rect 646 451 649 453
rect 651 451 654 453
rect 646 446 654 451
rect 646 444 649 446
rect 651 444 654 446
rect 646 442 654 444
rect 656 462 661 470
rect 668 468 675 470
rect 668 466 670 468
rect 672 466 675 468
rect 656 460 663 462
rect 656 458 659 460
rect 661 458 663 460
rect 656 453 663 458
rect 668 461 675 466
rect 668 459 670 461
rect 672 459 675 461
rect 668 457 675 459
rect 656 451 659 453
rect 661 451 663 453
rect 656 449 663 451
rect 656 442 661 449
rect 670 442 675 457
rect 677 453 685 470
rect 677 451 680 453
rect 682 451 685 453
rect 677 446 685 451
rect 677 444 680 446
rect 682 444 685 446
rect 677 442 685 444
rect 687 461 695 470
rect 687 459 690 461
rect 692 459 695 461
rect 687 454 695 459
rect 687 452 690 454
rect 692 452 695 454
rect 687 442 695 452
rect 697 453 713 470
rect 697 451 702 453
rect 704 451 713 453
rect 697 446 713 451
rect 697 444 702 446
rect 704 445 713 446
rect 715 445 720 470
rect 722 467 727 470
rect 722 465 730 467
rect 722 463 725 465
rect 727 463 730 465
rect 722 454 730 463
rect 732 454 743 467
rect 722 445 727 454
rect 734 446 743 454
rect 704 444 711 445
rect 697 442 711 444
rect 734 444 737 446
rect 739 444 743 446
rect 734 442 743 444
rect 745 465 752 467
rect 745 463 748 465
rect 750 463 752 465
rect 745 458 752 463
rect 745 456 748 458
rect 750 456 752 458
rect 745 454 752 456
rect 745 442 750 454
rect 82 431 89 433
rect 82 430 84 431
rect 73 424 78 430
rect 71 422 78 424
rect 71 420 73 422
rect 75 420 78 422
rect 71 415 78 420
rect 71 413 73 415
rect 75 413 78 415
rect 71 411 78 413
rect 73 402 78 411
rect 80 429 84 430
rect 86 430 89 431
rect 86 429 91 430
rect 80 402 91 429
rect 93 402 98 430
rect 100 424 105 430
rect 100 422 107 424
rect 100 420 103 422
rect 105 420 107 422
rect 100 418 107 420
rect 100 402 105 418
rect 114 415 119 430
rect 112 413 119 415
rect 112 411 114 413
rect 116 411 119 413
rect 112 406 119 411
rect 112 404 114 406
rect 116 404 119 406
rect 112 402 119 404
rect 121 428 129 430
rect 121 426 124 428
rect 126 426 129 428
rect 121 421 129 426
rect 121 419 124 421
rect 126 419 129 421
rect 121 402 129 419
rect 131 420 139 430
rect 131 418 134 420
rect 136 418 139 420
rect 131 413 139 418
rect 131 411 134 413
rect 136 411 139 413
rect 131 402 139 411
rect 141 428 155 430
rect 141 426 146 428
rect 148 427 155 428
rect 178 428 187 430
rect 148 426 157 427
rect 141 421 157 426
rect 141 419 146 421
rect 148 419 157 421
rect 141 402 157 419
rect 159 402 164 427
rect 166 418 171 427
rect 178 426 181 428
rect 183 426 187 428
rect 178 418 187 426
rect 166 409 174 418
rect 166 407 169 409
rect 171 407 174 409
rect 166 405 174 407
rect 176 405 187 418
rect 189 418 194 430
rect 189 416 196 418
rect 189 414 192 416
rect 194 414 196 416
rect 215 415 220 430
rect 189 409 196 414
rect 189 407 192 409
rect 194 407 196 409
rect 189 405 196 407
rect 213 413 220 415
rect 213 411 215 413
rect 217 411 220 413
rect 213 406 220 411
rect 166 402 171 405
rect 213 404 215 406
rect 217 404 220 406
rect 213 402 220 404
rect 222 428 230 430
rect 222 426 225 428
rect 227 426 230 428
rect 222 421 230 426
rect 222 419 225 421
rect 227 419 230 421
rect 222 402 230 419
rect 232 420 240 430
rect 232 418 235 420
rect 237 418 240 420
rect 232 413 240 418
rect 232 411 235 413
rect 237 411 240 413
rect 232 402 240 411
rect 242 428 256 430
rect 242 426 247 428
rect 249 427 256 428
rect 279 428 288 430
rect 249 426 258 427
rect 242 421 258 426
rect 242 419 247 421
rect 249 419 258 421
rect 242 402 258 419
rect 260 402 265 427
rect 267 418 272 427
rect 279 426 282 428
rect 284 426 288 428
rect 279 418 288 426
rect 267 409 275 418
rect 267 407 270 409
rect 272 407 275 409
rect 267 405 275 407
rect 277 405 288 418
rect 290 418 295 430
rect 290 416 297 418
rect 290 414 293 416
rect 295 414 297 416
rect 317 415 322 430
rect 290 409 297 414
rect 290 407 293 409
rect 295 407 297 409
rect 290 405 297 407
rect 315 413 322 415
rect 315 411 317 413
rect 319 411 322 413
rect 315 406 322 411
rect 267 402 272 405
rect 315 404 317 406
rect 319 404 322 406
rect 315 402 322 404
rect 324 428 332 430
rect 324 426 327 428
rect 329 426 332 428
rect 324 421 332 426
rect 324 419 327 421
rect 329 419 332 421
rect 324 402 332 419
rect 334 420 342 430
rect 334 418 337 420
rect 339 418 342 420
rect 334 413 342 418
rect 334 411 337 413
rect 339 411 342 413
rect 334 402 342 411
rect 344 428 358 430
rect 344 426 349 428
rect 351 427 358 428
rect 426 431 433 433
rect 426 430 428 431
rect 381 428 390 430
rect 351 426 360 427
rect 344 421 360 426
rect 344 419 349 421
rect 351 419 360 421
rect 344 402 360 419
rect 362 402 367 427
rect 369 418 374 427
rect 381 426 384 428
rect 386 426 390 428
rect 381 418 390 426
rect 369 409 377 418
rect 369 407 372 409
rect 374 407 377 409
rect 369 405 377 407
rect 379 405 390 418
rect 392 418 397 430
rect 417 424 422 430
rect 415 422 422 424
rect 415 420 417 422
rect 419 420 422 422
rect 392 416 399 418
rect 392 414 395 416
rect 397 414 399 416
rect 392 409 399 414
rect 415 415 422 420
rect 415 413 417 415
rect 419 413 422 415
rect 415 411 422 413
rect 392 407 395 409
rect 397 407 399 409
rect 392 405 399 407
rect 369 402 374 405
rect 417 402 422 411
rect 424 429 428 430
rect 430 430 433 431
rect 430 429 435 430
rect 424 402 435 429
rect 437 402 442 430
rect 444 424 449 430
rect 444 422 451 424
rect 444 420 447 422
rect 449 420 451 422
rect 444 418 451 420
rect 444 402 449 418
rect 470 415 475 430
rect 468 413 475 415
rect 468 411 470 413
rect 472 411 475 413
rect 468 406 475 411
rect 468 404 470 406
rect 472 404 475 406
rect 468 402 475 404
rect 477 428 485 430
rect 477 426 480 428
rect 482 426 485 428
rect 477 421 485 426
rect 477 419 480 421
rect 482 419 485 421
rect 477 402 485 419
rect 487 420 495 430
rect 487 418 490 420
rect 492 418 495 420
rect 487 413 495 418
rect 487 411 490 413
rect 492 411 495 413
rect 487 402 495 411
rect 497 428 511 430
rect 497 426 502 428
rect 504 427 511 428
rect 534 428 543 430
rect 504 426 513 427
rect 497 421 513 426
rect 497 419 502 421
rect 504 419 513 421
rect 497 402 513 419
rect 515 402 520 427
rect 522 418 527 427
rect 534 426 537 428
rect 539 426 543 428
rect 534 418 543 426
rect 522 409 530 418
rect 522 407 525 409
rect 527 407 530 409
rect 522 405 530 407
rect 532 405 543 418
rect 545 418 550 430
rect 545 416 552 418
rect 545 414 548 416
rect 550 414 552 416
rect 571 415 576 430
rect 545 409 552 414
rect 545 407 548 409
rect 550 407 552 409
rect 545 405 552 407
rect 569 413 576 415
rect 569 411 571 413
rect 573 411 576 413
rect 569 406 576 411
rect 522 402 527 405
rect 569 404 571 406
rect 573 404 576 406
rect 569 402 576 404
rect 578 428 586 430
rect 578 426 581 428
rect 583 426 586 428
rect 578 421 586 426
rect 578 419 581 421
rect 583 419 586 421
rect 578 402 586 419
rect 588 420 596 430
rect 588 418 591 420
rect 593 418 596 420
rect 588 413 596 418
rect 588 411 591 413
rect 593 411 596 413
rect 588 402 596 411
rect 598 428 612 430
rect 598 426 603 428
rect 605 427 612 428
rect 635 428 644 430
rect 605 426 614 427
rect 598 421 614 426
rect 598 419 603 421
rect 605 419 614 421
rect 598 402 614 419
rect 616 402 621 427
rect 623 418 628 427
rect 635 426 638 428
rect 640 426 644 428
rect 635 418 644 426
rect 623 409 631 418
rect 623 407 626 409
rect 628 407 631 409
rect 623 405 631 407
rect 633 405 644 418
rect 646 418 651 430
rect 646 416 653 418
rect 646 414 649 416
rect 651 414 653 416
rect 670 415 675 430
rect 646 409 653 414
rect 646 407 649 409
rect 651 407 653 409
rect 646 405 653 407
rect 668 413 675 415
rect 668 411 670 413
rect 672 411 675 413
rect 668 406 675 411
rect 623 402 628 405
rect 668 404 670 406
rect 672 404 675 406
rect 668 402 675 404
rect 677 428 685 430
rect 677 426 680 428
rect 682 426 685 428
rect 677 421 685 426
rect 677 419 680 421
rect 682 419 685 421
rect 677 402 685 419
rect 687 420 695 430
rect 687 418 690 420
rect 692 418 695 420
rect 687 413 695 418
rect 687 411 690 413
rect 692 411 695 413
rect 687 402 695 411
rect 697 428 711 430
rect 697 426 702 428
rect 704 427 711 428
rect 734 428 743 430
rect 704 426 713 427
rect 697 421 713 426
rect 697 419 702 421
rect 704 419 713 421
rect 697 402 713 419
rect 715 402 720 427
rect 722 418 727 427
rect 734 426 737 428
rect 739 426 743 428
rect 734 418 743 426
rect 722 409 730 418
rect 722 407 725 409
rect 727 407 730 409
rect 722 405 730 407
rect 732 405 743 418
rect 745 418 750 430
rect 745 416 752 418
rect 745 414 748 416
rect 750 414 752 416
rect 745 409 752 414
rect 745 407 748 409
rect 750 407 752 409
rect 745 405 752 407
rect 722 402 727 405
rect 73 324 80 326
rect 73 322 75 324
rect 77 322 80 324
rect 73 317 80 322
rect 73 315 75 317
rect 77 315 80 317
rect 73 313 80 315
rect 75 298 80 313
rect 82 309 90 326
rect 82 307 85 309
rect 87 307 90 309
rect 82 302 90 307
rect 82 300 85 302
rect 87 300 90 302
rect 82 298 90 300
rect 92 317 100 326
rect 92 315 95 317
rect 97 315 100 317
rect 92 310 100 315
rect 92 308 95 310
rect 97 308 100 310
rect 92 298 100 308
rect 102 309 118 326
rect 102 307 107 309
rect 109 307 118 309
rect 102 302 118 307
rect 102 300 107 302
rect 109 301 118 302
rect 120 301 125 326
rect 127 323 132 326
rect 127 321 135 323
rect 127 319 130 321
rect 132 319 135 321
rect 127 310 135 319
rect 137 310 148 323
rect 127 301 132 310
rect 139 302 148 310
rect 109 300 116 301
rect 102 298 116 300
rect 139 300 142 302
rect 144 300 148 302
rect 139 298 148 300
rect 150 321 157 323
rect 150 319 153 321
rect 155 319 157 321
rect 150 314 157 319
rect 163 317 168 326
rect 150 312 153 314
rect 155 312 157 314
rect 150 310 157 312
rect 161 315 168 317
rect 161 313 163 315
rect 165 313 168 315
rect 150 298 155 310
rect 161 308 168 313
rect 161 306 163 308
rect 165 306 168 308
rect 161 304 168 306
rect 163 298 168 304
rect 170 299 181 326
rect 170 298 174 299
rect 172 297 174 298
rect 176 298 181 299
rect 183 298 188 326
rect 190 310 195 326
rect 214 324 221 326
rect 214 322 216 324
rect 218 322 221 324
rect 214 317 221 322
rect 214 315 216 317
rect 218 315 221 317
rect 214 313 221 315
rect 190 308 197 310
rect 190 306 193 308
rect 195 306 197 308
rect 190 304 197 306
rect 190 298 195 304
rect 216 298 221 313
rect 223 309 231 326
rect 223 307 226 309
rect 228 307 231 309
rect 223 302 231 307
rect 223 300 226 302
rect 228 300 231 302
rect 223 298 231 300
rect 233 317 241 326
rect 233 315 236 317
rect 238 315 241 317
rect 233 310 241 315
rect 233 308 236 310
rect 238 308 241 310
rect 233 298 241 308
rect 243 309 259 326
rect 243 307 248 309
rect 250 307 259 309
rect 243 302 259 307
rect 243 300 248 302
rect 250 301 259 302
rect 261 301 266 326
rect 268 323 273 326
rect 339 323 344 326
rect 268 321 276 323
rect 268 319 271 321
rect 273 319 276 321
rect 268 310 276 319
rect 278 310 289 323
rect 268 301 273 310
rect 280 302 289 310
rect 250 300 257 301
rect 243 298 257 300
rect 176 297 179 298
rect 172 295 179 297
rect 280 300 283 302
rect 285 300 289 302
rect 280 298 289 300
rect 291 321 298 323
rect 291 319 294 321
rect 296 319 298 321
rect 291 314 298 319
rect 291 312 294 314
rect 296 312 298 314
rect 291 310 298 312
rect 314 321 321 323
rect 314 319 316 321
rect 318 319 321 321
rect 314 314 321 319
rect 314 312 316 314
rect 318 312 321 314
rect 314 310 321 312
rect 291 298 296 310
rect 316 298 321 310
rect 323 310 334 323
rect 336 321 344 323
rect 336 319 339 321
rect 341 319 344 321
rect 336 310 344 319
rect 323 302 332 310
rect 323 300 327 302
rect 329 300 332 302
rect 339 301 344 310
rect 346 301 351 326
rect 353 309 369 326
rect 353 307 362 309
rect 364 307 369 309
rect 353 302 369 307
rect 353 301 362 302
rect 323 298 332 300
rect 355 300 362 301
rect 364 300 369 302
rect 355 298 369 300
rect 371 317 379 326
rect 371 315 374 317
rect 376 315 379 317
rect 371 310 379 315
rect 371 308 374 310
rect 376 308 379 310
rect 371 298 379 308
rect 381 309 389 326
rect 381 307 384 309
rect 386 307 389 309
rect 381 302 389 307
rect 381 300 384 302
rect 386 300 389 302
rect 381 298 389 300
rect 391 324 398 326
rect 391 322 394 324
rect 396 322 398 324
rect 391 317 398 322
rect 417 317 422 326
rect 391 315 394 317
rect 396 315 398 317
rect 391 313 398 315
rect 415 315 422 317
rect 415 313 417 315
rect 419 313 422 315
rect 391 298 396 313
rect 415 308 422 313
rect 415 306 417 308
rect 419 306 422 308
rect 415 304 422 306
rect 417 298 422 304
rect 424 299 435 326
rect 424 298 428 299
rect 426 297 428 298
rect 430 298 435 299
rect 437 298 442 326
rect 444 310 449 326
rect 468 324 475 326
rect 468 322 470 324
rect 472 322 475 324
rect 468 317 475 322
rect 468 315 470 317
rect 472 315 475 317
rect 468 313 475 315
rect 444 308 451 310
rect 444 306 447 308
rect 449 306 451 308
rect 444 304 451 306
rect 444 298 449 304
rect 470 298 475 313
rect 477 309 485 326
rect 477 307 480 309
rect 482 307 485 309
rect 477 302 485 307
rect 477 300 480 302
rect 482 300 485 302
rect 477 298 485 300
rect 487 317 495 326
rect 487 315 490 317
rect 492 315 495 317
rect 487 310 495 315
rect 487 308 490 310
rect 492 308 495 310
rect 487 298 495 308
rect 497 309 513 326
rect 497 307 502 309
rect 504 307 513 309
rect 497 302 513 307
rect 497 300 502 302
rect 504 301 513 302
rect 515 301 520 326
rect 522 323 527 326
rect 569 324 576 326
rect 522 321 530 323
rect 522 319 525 321
rect 527 319 530 321
rect 522 310 530 319
rect 532 310 543 323
rect 522 301 527 310
rect 534 302 543 310
rect 504 300 511 301
rect 497 298 511 300
rect 430 297 433 298
rect 426 295 433 297
rect 534 300 537 302
rect 539 300 543 302
rect 534 298 543 300
rect 545 321 552 323
rect 545 319 548 321
rect 550 319 552 321
rect 545 314 552 319
rect 545 312 548 314
rect 550 312 552 314
rect 569 322 571 324
rect 573 322 576 324
rect 569 317 576 322
rect 569 315 571 317
rect 573 315 576 317
rect 569 313 576 315
rect 545 310 552 312
rect 545 298 550 310
rect 571 298 576 313
rect 578 309 586 326
rect 578 307 581 309
rect 583 307 586 309
rect 578 302 586 307
rect 578 300 581 302
rect 583 300 586 302
rect 578 298 586 300
rect 588 317 596 326
rect 588 315 591 317
rect 593 315 596 317
rect 588 310 596 315
rect 588 308 591 310
rect 593 308 596 310
rect 588 298 596 308
rect 598 309 614 326
rect 598 307 603 309
rect 605 307 614 309
rect 598 302 614 307
rect 598 300 603 302
rect 605 301 614 302
rect 616 301 621 326
rect 623 323 628 326
rect 668 324 675 326
rect 623 321 631 323
rect 623 319 626 321
rect 628 319 631 321
rect 623 310 631 319
rect 633 310 644 323
rect 623 301 628 310
rect 635 302 644 310
rect 605 300 612 301
rect 598 298 612 300
rect 635 300 638 302
rect 640 300 644 302
rect 635 298 644 300
rect 646 321 653 323
rect 646 319 649 321
rect 651 319 653 321
rect 646 314 653 319
rect 646 312 649 314
rect 651 312 653 314
rect 668 322 670 324
rect 672 322 675 324
rect 668 317 675 322
rect 668 315 670 317
rect 672 315 675 317
rect 668 313 675 315
rect 646 310 653 312
rect 646 298 651 310
rect 670 298 675 313
rect 677 309 685 326
rect 677 307 680 309
rect 682 307 685 309
rect 677 302 685 307
rect 677 300 680 302
rect 682 300 685 302
rect 677 298 685 300
rect 687 317 695 326
rect 687 315 690 317
rect 692 315 695 317
rect 687 310 695 315
rect 687 308 690 310
rect 692 308 695 310
rect 687 298 695 308
rect 697 309 713 326
rect 697 307 702 309
rect 704 307 713 309
rect 697 302 713 307
rect 697 300 702 302
rect 704 301 713 302
rect 715 301 720 326
rect 722 323 727 326
rect 722 321 730 323
rect 722 319 725 321
rect 727 319 730 321
rect 722 310 730 319
rect 732 310 743 323
rect 722 301 727 310
rect 734 302 743 310
rect 704 300 711 301
rect 697 298 711 300
rect 734 300 737 302
rect 739 300 743 302
rect 734 298 743 300
rect 745 321 752 323
rect 745 319 748 321
rect 750 319 752 321
rect 745 314 752 319
rect 745 312 748 314
rect 750 312 752 314
rect 745 310 752 312
rect 745 298 750 310
rect 82 287 89 289
rect 82 286 84 287
rect 73 280 78 286
rect 71 278 78 280
rect 71 276 73 278
rect 75 276 78 278
rect 71 271 78 276
rect 71 269 73 271
rect 75 269 78 271
rect 71 267 78 269
rect 73 258 78 267
rect 80 285 84 286
rect 86 286 89 287
rect 86 285 91 286
rect 80 258 91 285
rect 93 258 98 286
rect 100 280 105 286
rect 100 278 107 280
rect 100 276 103 278
rect 105 276 107 278
rect 100 274 107 276
rect 100 258 105 274
rect 114 271 119 286
rect 112 269 119 271
rect 112 267 114 269
rect 116 267 119 269
rect 112 262 119 267
rect 112 260 114 262
rect 116 260 119 262
rect 112 258 119 260
rect 121 284 129 286
rect 121 282 124 284
rect 126 282 129 284
rect 121 277 129 282
rect 121 275 124 277
rect 126 275 129 277
rect 121 258 129 275
rect 131 276 139 286
rect 131 274 134 276
rect 136 274 139 276
rect 131 269 139 274
rect 131 267 134 269
rect 136 267 139 269
rect 131 258 139 267
rect 141 284 155 286
rect 141 282 146 284
rect 148 283 155 284
rect 178 284 187 286
rect 148 282 157 283
rect 141 277 157 282
rect 141 275 146 277
rect 148 275 157 277
rect 141 258 157 275
rect 159 258 164 283
rect 166 274 171 283
rect 178 282 181 284
rect 183 282 187 284
rect 178 274 187 282
rect 166 265 174 274
rect 166 263 169 265
rect 171 263 174 265
rect 166 261 174 263
rect 176 261 187 274
rect 189 274 194 286
rect 189 272 196 274
rect 189 270 192 272
rect 194 270 196 272
rect 215 271 220 286
rect 189 265 196 270
rect 189 263 192 265
rect 194 263 196 265
rect 189 261 196 263
rect 213 269 220 271
rect 213 267 215 269
rect 217 267 220 269
rect 213 262 220 267
rect 166 258 171 261
rect 213 260 215 262
rect 217 260 220 262
rect 213 258 220 260
rect 222 284 230 286
rect 222 282 225 284
rect 227 282 230 284
rect 222 277 230 282
rect 222 275 225 277
rect 227 275 230 277
rect 222 258 230 275
rect 232 276 240 286
rect 232 274 235 276
rect 237 274 240 276
rect 232 269 240 274
rect 232 267 235 269
rect 237 267 240 269
rect 232 258 240 267
rect 242 284 256 286
rect 242 282 247 284
rect 249 283 256 284
rect 279 284 288 286
rect 249 282 258 283
rect 242 277 258 282
rect 242 275 247 277
rect 249 275 258 277
rect 242 258 258 275
rect 260 258 265 283
rect 267 274 272 283
rect 279 282 282 284
rect 284 282 288 284
rect 279 274 288 282
rect 267 265 275 274
rect 267 263 270 265
rect 272 263 275 265
rect 267 261 275 263
rect 277 261 288 274
rect 290 274 295 286
rect 290 272 297 274
rect 290 270 293 272
rect 295 270 297 272
rect 316 271 321 286
rect 290 265 297 270
rect 290 263 293 265
rect 295 263 297 265
rect 290 261 297 263
rect 314 269 321 271
rect 314 267 316 269
rect 318 267 321 269
rect 314 262 321 267
rect 267 258 272 261
rect 314 260 316 262
rect 318 260 321 262
rect 314 258 321 260
rect 323 284 331 286
rect 323 282 326 284
rect 328 282 331 284
rect 323 277 331 282
rect 323 275 326 277
rect 328 275 331 277
rect 323 258 331 275
rect 333 276 341 286
rect 333 274 336 276
rect 338 274 341 276
rect 333 269 341 274
rect 333 267 336 269
rect 338 267 341 269
rect 333 258 341 267
rect 343 284 357 286
rect 343 282 348 284
rect 350 283 357 284
rect 425 287 432 289
rect 425 286 427 287
rect 380 284 389 286
rect 350 282 359 283
rect 343 277 359 282
rect 343 275 348 277
rect 350 275 359 277
rect 343 258 359 275
rect 361 258 366 283
rect 368 274 373 283
rect 380 282 383 284
rect 385 282 389 284
rect 380 274 389 282
rect 368 265 376 274
rect 368 263 371 265
rect 373 263 376 265
rect 368 261 376 263
rect 378 261 389 274
rect 391 274 396 286
rect 416 280 421 286
rect 414 278 421 280
rect 414 276 416 278
rect 418 276 421 278
rect 391 272 398 274
rect 391 270 394 272
rect 396 270 398 272
rect 391 265 398 270
rect 414 271 421 276
rect 414 269 416 271
rect 418 269 421 271
rect 414 267 421 269
rect 391 263 394 265
rect 396 263 398 265
rect 391 261 398 263
rect 368 258 373 261
rect 416 258 421 267
rect 423 285 427 286
rect 429 286 432 287
rect 429 285 434 286
rect 423 258 434 285
rect 436 258 441 286
rect 443 280 448 286
rect 443 278 450 280
rect 443 276 446 278
rect 448 276 450 278
rect 443 274 450 276
rect 443 258 448 274
rect 469 271 474 286
rect 467 269 474 271
rect 467 267 469 269
rect 471 267 474 269
rect 467 262 474 267
rect 467 260 469 262
rect 471 260 474 262
rect 467 258 474 260
rect 476 284 484 286
rect 476 282 479 284
rect 481 282 484 284
rect 476 277 484 282
rect 476 275 479 277
rect 481 275 484 277
rect 476 258 484 275
rect 486 276 494 286
rect 486 274 489 276
rect 491 274 494 276
rect 486 269 494 274
rect 486 267 489 269
rect 491 267 494 269
rect 486 258 494 267
rect 496 284 510 286
rect 496 282 501 284
rect 503 283 510 284
rect 533 284 542 286
rect 503 282 512 283
rect 496 277 512 282
rect 496 275 501 277
rect 503 275 512 277
rect 496 258 512 275
rect 514 258 519 283
rect 521 274 526 283
rect 533 282 536 284
rect 538 282 542 284
rect 533 274 542 282
rect 521 265 529 274
rect 521 263 524 265
rect 526 263 529 265
rect 521 261 529 263
rect 531 261 542 274
rect 544 274 549 286
rect 544 272 551 274
rect 544 270 547 272
rect 549 270 551 272
rect 570 271 575 286
rect 544 265 551 270
rect 544 263 547 265
rect 549 263 551 265
rect 544 261 551 263
rect 568 269 575 271
rect 568 267 570 269
rect 572 267 575 269
rect 568 262 575 267
rect 521 258 526 261
rect 568 260 570 262
rect 572 260 575 262
rect 568 258 575 260
rect 577 284 585 286
rect 577 282 580 284
rect 582 282 585 284
rect 577 277 585 282
rect 577 275 580 277
rect 582 275 585 277
rect 577 258 585 275
rect 587 276 595 286
rect 587 274 590 276
rect 592 274 595 276
rect 587 269 595 274
rect 587 267 590 269
rect 592 267 595 269
rect 587 258 595 267
rect 597 284 611 286
rect 597 282 602 284
rect 604 283 611 284
rect 634 284 643 286
rect 604 282 613 283
rect 597 277 613 282
rect 597 275 602 277
rect 604 275 613 277
rect 597 258 613 275
rect 615 258 620 283
rect 622 274 627 283
rect 634 282 637 284
rect 639 282 643 284
rect 634 274 643 282
rect 622 265 630 274
rect 622 263 625 265
rect 627 263 630 265
rect 622 261 630 263
rect 632 261 643 274
rect 645 274 650 286
rect 645 272 652 274
rect 645 270 648 272
rect 650 270 652 272
rect 669 271 674 286
rect 645 265 652 270
rect 645 263 648 265
rect 650 263 652 265
rect 645 261 652 263
rect 667 269 674 271
rect 667 267 669 269
rect 671 267 674 269
rect 667 262 674 267
rect 622 258 627 261
rect 667 260 669 262
rect 671 260 674 262
rect 667 258 674 260
rect 676 284 684 286
rect 676 282 679 284
rect 681 282 684 284
rect 676 277 684 282
rect 676 275 679 277
rect 681 275 684 277
rect 676 258 684 275
rect 686 276 694 286
rect 686 274 689 276
rect 691 274 694 276
rect 686 269 694 274
rect 686 267 689 269
rect 691 267 694 269
rect 686 258 694 267
rect 696 284 710 286
rect 696 282 701 284
rect 703 283 710 284
rect 733 284 742 286
rect 703 282 712 283
rect 696 277 712 282
rect 696 275 701 277
rect 703 275 712 277
rect 696 258 712 275
rect 714 258 719 283
rect 721 274 726 283
rect 733 282 736 284
rect 738 282 742 284
rect 733 274 742 282
rect 721 265 729 274
rect 721 263 724 265
rect 726 263 729 265
rect 721 261 729 263
rect 731 261 742 274
rect 744 274 749 286
rect 744 272 751 274
rect 744 270 747 272
rect 749 270 751 272
rect 744 265 751 270
rect 744 263 747 265
rect 749 263 751 265
rect 744 261 751 263
rect 721 258 726 261
<< alu1 >>
rect 402 581 406 582
rect 402 580 403 581
rect 67 579 403 580
rect 405 580 406 581
rect 448 581 452 582
rect 448 580 449 581
rect 405 579 449 580
rect 451 580 452 581
rect 493 581 497 582
rect 493 580 494 581
rect 451 579 494 580
rect 496 580 497 581
rect 566 581 570 582
rect 566 580 567 581
rect 496 579 567 580
rect 569 580 570 581
rect 569 579 756 580
rect 67 578 756 579
rect 67 577 108 578
rect 67 575 68 577
rect 70 576 108 577
rect 110 577 753 578
rect 110 576 146 577
rect 70 575 146 576
rect 148 575 217 577
rect 219 575 282 577
rect 284 575 335 577
rect 337 575 370 577
rect 372 575 632 577
rect 634 576 753 577
rect 755 576 756 578
rect 634 575 756 576
rect 67 572 756 575
rect 102 565 107 567
rect 102 563 103 565
rect 105 563 107 565
rect 71 550 75 559
rect 102 558 107 563
rect 142 565 147 567
rect 142 563 143 565
rect 145 563 147 565
rect 102 556 103 558
rect 105 556 107 558
rect 102 554 107 556
rect 71 549 84 550
rect 71 547 76 549
rect 78 547 81 549
rect 83 547 84 549
rect 71 546 84 547
rect 78 541 92 542
rect 78 539 86 541
rect 88 539 92 541
rect 78 538 92 539
rect 78 532 83 538
rect 78 530 79 532
rect 81 530 83 532
rect 78 529 83 530
rect 103 532 107 554
rect 111 550 115 559
rect 142 558 147 563
rect 223 562 236 566
rect 142 556 143 558
rect 145 556 147 558
rect 142 554 147 556
rect 111 549 124 550
rect 111 547 112 549
rect 114 547 116 549
rect 118 547 124 549
rect 111 546 124 547
rect 105 530 107 532
rect 103 527 107 530
rect 118 541 132 542
rect 118 539 126 541
rect 128 539 132 541
rect 118 538 132 539
rect 118 532 123 538
rect 118 530 119 532
rect 121 530 123 532
rect 118 529 123 530
rect 95 524 107 527
rect 143 532 147 554
rect 145 530 147 532
rect 143 527 147 530
rect 95 522 103 524
rect 105 522 107 524
rect 135 524 147 527
rect 135 522 143 524
rect 145 522 147 524
rect 151 557 157 559
rect 231 560 236 562
rect 231 558 232 560
rect 234 558 236 560
rect 151 555 154 557
rect 156 555 157 557
rect 151 550 157 555
rect 151 548 154 550
rect 156 548 157 550
rect 151 546 157 548
rect 151 526 155 546
rect 167 549 205 550
rect 167 547 168 549
rect 170 547 205 549
rect 167 546 205 547
rect 200 543 205 546
rect 175 541 190 542
rect 175 539 179 541
rect 181 539 186 541
rect 188 539 190 541
rect 175 538 190 539
rect 200 541 208 543
rect 200 539 205 541
rect 207 539 208 541
rect 184 532 188 538
rect 200 537 208 539
rect 231 553 236 558
rect 231 551 232 553
rect 234 551 236 553
rect 231 549 236 551
rect 184 530 185 532
rect 187 530 188 532
rect 184 529 188 530
rect 151 525 173 526
rect 151 523 154 525
rect 156 523 170 525
rect 172 523 173 525
rect 151 522 173 523
rect 232 527 236 549
rect 231 525 236 527
rect 231 523 232 525
rect 234 523 236 525
rect 95 521 107 522
rect 135 521 147 522
rect 231 521 236 523
rect 248 562 261 566
rect 337 565 342 567
rect 337 563 339 565
rect 341 563 342 565
rect 248 560 253 562
rect 248 558 250 560
rect 252 558 253 560
rect 248 553 253 558
rect 248 551 250 553
rect 252 551 253 553
rect 248 549 253 551
rect 248 527 252 549
rect 279 549 317 550
rect 279 547 314 549
rect 316 547 317 549
rect 279 546 317 547
rect 279 543 284 546
rect 276 541 284 543
rect 276 539 277 541
rect 279 539 284 541
rect 276 537 284 539
rect 294 541 309 542
rect 294 539 296 541
rect 298 539 303 541
rect 305 539 309 541
rect 294 538 309 539
rect 248 525 253 527
rect 296 532 300 538
rect 327 557 333 559
rect 327 555 328 557
rect 330 555 333 557
rect 327 550 333 555
rect 327 548 328 550
rect 330 548 333 550
rect 327 546 333 548
rect 296 530 297 532
rect 299 530 300 532
rect 296 529 300 530
rect 329 526 333 546
rect 248 523 250 525
rect 252 523 253 525
rect 248 521 253 523
rect 311 525 333 526
rect 311 523 312 525
rect 314 523 328 525
rect 330 523 333 525
rect 311 522 333 523
rect 337 558 342 563
rect 377 565 382 567
rect 377 563 379 565
rect 381 563 382 565
rect 337 556 339 558
rect 341 556 342 558
rect 337 554 342 556
rect 337 532 341 554
rect 369 550 373 559
rect 360 549 373 550
rect 360 547 366 549
rect 368 547 370 549
rect 372 547 373 549
rect 360 546 373 547
rect 377 558 382 563
rect 418 562 431 566
rect 507 565 512 567
rect 507 563 509 565
rect 511 563 512 565
rect 418 560 423 562
rect 377 556 379 558
rect 381 556 382 558
rect 377 554 382 556
rect 352 541 366 542
rect 352 539 356 541
rect 358 539 366 541
rect 352 538 366 539
rect 337 530 339 532
rect 337 527 341 530
rect 337 524 349 527
rect 337 522 339 524
rect 341 522 349 524
rect 361 532 366 538
rect 361 530 363 532
rect 365 530 366 532
rect 361 529 366 530
rect 377 532 381 554
rect 409 550 413 559
rect 400 549 413 550
rect 400 547 401 549
rect 403 547 406 549
rect 408 547 413 549
rect 400 546 413 547
rect 418 558 420 560
rect 422 558 423 560
rect 418 553 423 558
rect 418 551 420 553
rect 422 551 423 553
rect 418 549 423 551
rect 392 541 406 542
rect 392 539 396 541
rect 398 539 406 541
rect 392 538 406 539
rect 377 530 379 532
rect 377 527 381 530
rect 377 524 389 527
rect 377 522 379 524
rect 381 522 389 524
rect 401 532 406 538
rect 401 530 403 532
rect 405 530 406 532
rect 401 529 406 530
rect 418 527 422 549
rect 449 549 487 550
rect 449 547 484 549
rect 486 547 487 549
rect 449 546 487 547
rect 449 543 454 546
rect 446 541 454 543
rect 446 539 447 541
rect 449 539 454 541
rect 446 537 454 539
rect 464 541 479 542
rect 464 539 466 541
rect 468 539 473 541
rect 475 539 479 541
rect 464 538 479 539
rect 418 525 423 527
rect 466 532 470 538
rect 497 557 503 559
rect 497 555 498 557
rect 500 555 503 557
rect 497 550 503 555
rect 497 548 498 550
rect 500 548 503 550
rect 497 546 503 548
rect 466 530 467 532
rect 469 530 470 532
rect 466 529 470 530
rect 499 526 503 546
rect 418 523 420 525
rect 422 523 423 525
rect 337 521 349 522
rect 377 521 389 522
rect 418 521 423 523
rect 481 525 503 526
rect 481 523 482 525
rect 484 523 498 525
rect 500 523 503 525
rect 481 522 503 523
rect 507 558 512 563
rect 547 565 552 567
rect 547 563 549 565
rect 551 563 552 565
rect 507 556 509 558
rect 511 556 512 558
rect 507 554 512 556
rect 507 532 511 554
rect 539 550 543 559
rect 530 549 543 550
rect 530 547 536 549
rect 538 547 540 549
rect 542 547 543 549
rect 530 546 543 547
rect 547 558 552 563
rect 618 565 623 567
rect 618 563 619 565
rect 621 563 623 565
rect 547 556 549 558
rect 551 556 552 558
rect 547 554 552 556
rect 522 541 536 542
rect 522 539 526 541
rect 528 539 536 541
rect 522 538 536 539
rect 507 530 509 532
rect 507 527 511 530
rect 507 524 519 527
rect 507 522 509 524
rect 511 522 519 524
rect 531 532 536 538
rect 531 530 533 532
rect 535 530 536 532
rect 531 529 536 530
rect 547 532 551 554
rect 579 550 583 559
rect 570 549 583 550
rect 570 547 571 549
rect 573 547 576 549
rect 578 547 583 549
rect 570 546 583 547
rect 587 550 591 559
rect 618 558 623 563
rect 658 565 663 567
rect 658 563 659 565
rect 661 563 663 565
rect 618 556 619 558
rect 621 556 623 558
rect 618 554 623 556
rect 587 549 600 550
rect 587 547 592 549
rect 594 547 597 549
rect 599 547 600 549
rect 587 546 600 547
rect 562 541 576 542
rect 562 539 566 541
rect 568 539 576 541
rect 562 538 576 539
rect 547 530 549 532
rect 547 527 551 530
rect 547 524 559 527
rect 547 522 549 524
rect 551 522 559 524
rect 571 532 576 538
rect 571 530 573 532
rect 575 530 576 532
rect 571 529 576 530
rect 594 541 608 542
rect 594 539 602 541
rect 604 539 608 541
rect 594 538 608 539
rect 594 532 599 538
rect 594 530 595 532
rect 597 530 599 532
rect 594 529 599 530
rect 619 532 623 554
rect 627 550 631 559
rect 658 558 663 563
rect 739 562 752 566
rect 658 556 659 558
rect 661 556 663 558
rect 658 554 663 556
rect 627 549 640 550
rect 627 547 628 549
rect 630 547 632 549
rect 634 547 640 549
rect 627 546 640 547
rect 621 530 623 532
rect 619 527 623 530
rect 634 541 648 542
rect 634 539 642 541
rect 644 539 648 541
rect 634 538 648 539
rect 634 532 639 538
rect 634 530 635 532
rect 637 530 639 532
rect 634 529 639 530
rect 611 524 623 527
rect 659 532 663 554
rect 661 530 663 532
rect 659 527 663 530
rect 611 522 619 524
rect 621 522 623 524
rect 651 524 663 527
rect 651 522 659 524
rect 661 522 663 524
rect 667 557 673 559
rect 747 560 752 562
rect 747 558 748 560
rect 750 558 752 560
rect 667 555 670 557
rect 672 555 673 557
rect 667 550 673 555
rect 667 548 670 550
rect 672 548 673 550
rect 667 546 673 548
rect 667 526 671 546
rect 683 549 721 550
rect 683 547 684 549
rect 686 547 721 549
rect 683 546 721 547
rect 716 543 721 546
rect 691 541 706 542
rect 691 539 695 541
rect 697 539 702 541
rect 704 539 706 541
rect 691 538 706 539
rect 716 541 724 543
rect 716 539 721 541
rect 723 539 724 541
rect 700 532 704 538
rect 716 537 724 539
rect 747 553 752 558
rect 747 551 748 553
rect 750 551 752 553
rect 747 549 752 551
rect 700 530 701 532
rect 703 530 704 532
rect 700 529 704 530
rect 667 525 689 526
rect 667 523 670 525
rect 672 523 686 525
rect 688 523 689 525
rect 667 522 689 523
rect 748 527 752 549
rect 747 525 752 527
rect 747 523 748 525
rect 750 523 752 525
rect 507 521 519 522
rect 547 521 559 522
rect 611 521 623 522
rect 651 521 663 522
rect 747 521 752 523
rect 67 515 756 516
rect 67 513 92 515
rect 94 513 132 515
rect 134 513 350 515
rect 352 513 390 515
rect 392 513 520 515
rect 522 513 560 515
rect 562 513 608 515
rect 610 513 648 515
rect 650 513 756 515
rect 67 509 756 513
rect 67 507 68 509
rect 70 507 129 509
rect 131 507 193 509
rect 195 507 257 509
rect 259 507 320 509
rect 322 507 355 509
rect 357 507 387 509
rect 389 507 428 509
rect 430 507 459 509
rect 461 507 516 509
rect 518 507 606 509
rect 608 507 709 509
rect 711 507 753 509
rect 755 507 756 509
rect 67 503 756 507
rect 67 501 92 503
rect 94 501 132 503
rect 134 501 350 503
rect 352 501 390 503
rect 392 501 520 503
rect 522 501 560 503
rect 562 501 608 503
rect 610 501 648 503
rect 650 501 756 503
rect 67 500 756 501
rect 95 494 107 495
rect 135 494 147 495
rect 78 486 83 487
rect 78 484 79 486
rect 81 484 83 486
rect 78 478 83 484
rect 95 492 103 494
rect 105 492 107 494
rect 95 489 107 492
rect 103 486 107 489
rect 105 484 107 486
rect 78 477 92 478
rect 78 475 86 477
rect 88 475 92 477
rect 78 474 92 475
rect 71 469 84 470
rect 71 467 76 469
rect 78 467 81 469
rect 83 467 84 469
rect 71 466 84 467
rect 103 477 107 484
rect 103 475 104 477
rect 106 475 107 477
rect 71 457 75 466
rect 103 462 107 475
rect 118 486 123 487
rect 118 484 119 486
rect 121 484 123 486
rect 118 478 123 484
rect 135 492 143 494
rect 145 492 147 494
rect 135 489 147 492
rect 143 486 147 489
rect 145 484 147 486
rect 118 477 132 478
rect 118 475 126 477
rect 128 475 132 477
rect 118 474 132 475
rect 102 460 107 462
rect 102 458 103 460
rect 105 458 107 460
rect 102 453 107 458
rect 111 469 124 470
rect 111 467 112 469
rect 114 467 116 469
rect 118 467 124 469
rect 111 466 124 467
rect 111 457 115 466
rect 143 462 147 484
rect 142 460 147 462
rect 142 458 143 460
rect 145 458 147 460
rect 102 451 103 453
rect 105 451 107 453
rect 102 449 107 451
rect 142 453 147 458
rect 151 493 173 494
rect 151 491 154 493
rect 156 491 173 493
rect 151 490 173 491
rect 231 493 236 495
rect 231 491 232 493
rect 234 491 236 493
rect 151 470 155 490
rect 151 468 157 470
rect 151 466 154 468
rect 156 466 157 468
rect 151 461 157 466
rect 151 459 154 461
rect 156 459 157 461
rect 151 457 157 459
rect 184 478 188 487
rect 231 489 236 491
rect 175 477 190 478
rect 175 475 176 477
rect 178 475 179 477
rect 181 475 186 477
rect 188 475 190 477
rect 175 474 190 475
rect 200 477 208 479
rect 200 475 205 477
rect 207 475 208 477
rect 200 473 208 475
rect 200 470 205 473
rect 167 469 205 470
rect 167 467 168 469
rect 170 467 205 469
rect 167 466 205 467
rect 232 467 236 489
rect 231 465 236 467
rect 231 463 232 465
rect 234 463 236 465
rect 231 458 236 463
rect 231 456 232 458
rect 234 456 236 458
rect 231 454 236 456
rect 142 451 143 453
rect 145 451 147 453
rect 142 449 147 451
rect 223 450 236 454
rect 248 493 253 495
rect 337 494 349 495
rect 377 494 389 495
rect 248 491 250 493
rect 252 491 253 493
rect 248 489 253 491
rect 248 467 252 489
rect 311 493 333 494
rect 311 491 328 493
rect 330 491 333 493
rect 311 490 333 491
rect 248 465 253 467
rect 248 463 250 465
rect 252 463 253 465
rect 248 458 253 463
rect 276 477 284 479
rect 296 478 300 487
rect 276 475 277 477
rect 279 475 284 477
rect 276 473 284 475
rect 294 477 309 478
rect 294 475 296 477
rect 298 475 303 477
rect 305 475 306 477
rect 308 475 309 477
rect 294 474 309 475
rect 279 470 284 473
rect 279 469 317 470
rect 279 467 314 469
rect 316 467 317 469
rect 279 466 317 467
rect 329 470 333 490
rect 327 468 333 470
rect 327 466 328 468
rect 330 466 333 468
rect 327 461 333 466
rect 327 459 328 461
rect 330 459 333 461
rect 248 456 250 458
rect 252 456 253 458
rect 248 454 253 456
rect 327 457 333 459
rect 337 492 339 494
rect 341 492 349 494
rect 337 489 349 492
rect 377 492 379 494
rect 381 492 389 494
rect 337 486 341 489
rect 337 484 339 486
rect 337 462 341 484
rect 377 489 389 492
rect 418 493 423 495
rect 507 494 519 495
rect 547 494 559 495
rect 611 494 623 495
rect 651 494 663 495
rect 418 491 420 493
rect 422 491 423 493
rect 361 486 366 487
rect 361 484 363 486
rect 365 484 366 486
rect 361 478 366 484
rect 352 477 366 478
rect 352 475 356 477
rect 358 475 366 477
rect 352 474 366 475
rect 377 486 381 489
rect 377 484 379 486
rect 360 469 373 470
rect 360 467 366 469
rect 368 467 370 469
rect 372 467 373 469
rect 360 466 373 467
rect 337 460 342 462
rect 337 458 339 460
rect 341 458 342 460
rect 248 450 261 454
rect 337 453 342 458
rect 369 457 373 466
rect 377 462 381 484
rect 418 489 423 491
rect 401 486 406 487
rect 401 484 403 486
rect 405 484 406 486
rect 401 478 406 484
rect 392 477 406 478
rect 392 475 396 477
rect 398 475 406 477
rect 392 474 406 475
rect 400 469 413 470
rect 400 467 401 469
rect 403 467 406 469
rect 408 467 413 469
rect 400 466 413 467
rect 377 460 382 462
rect 377 458 379 460
rect 381 458 382 460
rect 337 451 339 453
rect 341 451 342 453
rect 337 449 342 451
rect 377 456 382 458
rect 377 454 379 456
rect 381 454 382 456
rect 409 457 413 466
rect 418 467 422 489
rect 481 493 503 494
rect 481 491 498 493
rect 500 491 503 493
rect 481 490 503 491
rect 418 465 423 467
rect 418 463 420 465
rect 422 463 423 465
rect 418 458 423 463
rect 446 477 454 479
rect 466 478 470 487
rect 499 485 503 490
rect 499 483 500 485
rect 502 483 503 485
rect 446 475 447 477
rect 449 475 454 477
rect 446 473 454 475
rect 464 477 479 478
rect 464 475 466 477
rect 468 475 473 477
rect 475 475 476 477
rect 478 475 479 477
rect 464 474 479 475
rect 449 470 454 473
rect 449 469 487 470
rect 449 467 484 469
rect 486 467 487 469
rect 449 466 487 467
rect 499 470 503 483
rect 497 468 503 470
rect 497 466 498 468
rect 500 466 503 468
rect 497 461 503 466
rect 497 459 498 461
rect 500 459 503 461
rect 377 453 382 454
rect 377 451 379 453
rect 381 451 382 453
rect 377 449 382 451
rect 418 456 420 458
rect 422 456 423 458
rect 418 454 423 456
rect 497 457 503 459
rect 507 492 509 494
rect 511 492 519 494
rect 507 489 519 492
rect 547 492 549 494
rect 551 492 559 494
rect 507 486 511 489
rect 507 484 509 486
rect 507 462 511 484
rect 547 489 559 492
rect 531 486 536 487
rect 531 484 533 486
rect 535 484 536 486
rect 531 478 536 484
rect 522 477 536 478
rect 522 475 526 477
rect 528 475 536 477
rect 522 474 536 475
rect 547 486 551 489
rect 547 484 549 486
rect 547 477 551 484
rect 571 486 576 487
rect 571 484 573 486
rect 575 484 576 486
rect 547 475 548 477
rect 550 475 551 477
rect 530 469 543 470
rect 530 467 536 469
rect 538 467 540 469
rect 542 467 543 469
rect 530 466 543 467
rect 507 460 512 462
rect 507 458 509 460
rect 511 458 512 460
rect 418 450 431 454
rect 507 453 512 458
rect 539 457 543 466
rect 547 462 551 475
rect 571 478 576 484
rect 562 477 576 478
rect 562 475 566 477
rect 568 475 576 477
rect 562 474 576 475
rect 594 486 599 487
rect 594 484 595 486
rect 597 484 599 486
rect 594 478 599 484
rect 611 492 619 494
rect 621 492 623 494
rect 611 489 623 492
rect 619 486 623 489
rect 621 484 623 486
rect 594 477 608 478
rect 594 475 602 477
rect 604 475 608 477
rect 594 474 608 475
rect 570 469 583 470
rect 570 467 571 469
rect 573 467 576 469
rect 578 467 583 469
rect 570 466 583 467
rect 547 460 552 462
rect 547 458 549 460
rect 551 458 552 460
rect 507 451 509 453
rect 511 451 512 453
rect 507 449 512 451
rect 547 453 552 458
rect 579 457 583 466
rect 587 469 600 470
rect 587 467 592 469
rect 594 467 597 469
rect 599 467 600 469
rect 587 466 600 467
rect 587 457 591 466
rect 619 462 623 484
rect 634 486 639 487
rect 634 484 635 486
rect 637 484 639 486
rect 634 478 639 484
rect 651 492 659 494
rect 661 492 663 494
rect 651 489 663 492
rect 659 486 663 489
rect 661 484 663 486
rect 634 477 648 478
rect 634 475 642 477
rect 644 475 648 477
rect 634 474 648 475
rect 618 460 623 462
rect 618 458 619 460
rect 621 458 623 460
rect 547 451 549 453
rect 551 451 552 453
rect 547 449 552 451
rect 618 453 623 458
rect 627 469 640 470
rect 627 467 628 469
rect 630 467 632 469
rect 634 467 640 469
rect 627 466 640 467
rect 627 457 631 466
rect 659 462 663 484
rect 658 460 663 462
rect 658 458 659 460
rect 661 458 663 460
rect 618 451 619 453
rect 621 451 623 453
rect 618 449 623 451
rect 658 453 663 458
rect 667 493 689 494
rect 667 491 670 493
rect 672 491 689 493
rect 667 490 689 491
rect 747 493 752 495
rect 747 491 748 493
rect 750 491 752 493
rect 667 470 671 490
rect 667 468 673 470
rect 667 466 670 468
rect 672 466 673 468
rect 667 461 673 466
rect 667 459 670 461
rect 672 459 673 461
rect 667 457 673 459
rect 700 478 704 487
rect 747 489 752 491
rect 691 477 706 478
rect 691 475 692 477
rect 694 475 695 477
rect 697 475 702 477
rect 704 475 706 477
rect 691 474 706 475
rect 716 477 724 479
rect 716 475 721 477
rect 723 475 724 477
rect 716 473 724 475
rect 716 470 721 473
rect 683 469 721 470
rect 683 467 684 469
rect 686 467 721 469
rect 683 466 721 467
rect 748 467 752 489
rect 747 465 752 467
rect 747 463 748 465
rect 750 463 752 465
rect 747 458 752 463
rect 747 456 748 458
rect 750 456 752 458
rect 747 454 752 456
rect 658 451 659 453
rect 661 451 663 453
rect 658 449 663 451
rect 739 453 752 454
rect 739 451 740 453
rect 742 451 752 453
rect 739 450 752 451
rect 67 438 756 444
rect 67 437 753 438
rect 67 436 108 437
rect 67 434 68 436
rect 70 435 108 436
rect 110 435 146 437
rect 148 435 217 437
rect 219 435 282 437
rect 284 435 335 437
rect 337 436 449 437
rect 337 435 370 436
rect 70 434 370 435
rect 372 434 402 436
rect 404 435 449 436
rect 451 435 494 437
rect 496 436 753 437
rect 755 436 756 438
rect 496 435 567 436
rect 404 434 567 435
rect 569 434 632 436
rect 634 434 756 436
rect 67 431 756 434
rect 67 429 84 431
rect 86 429 428 431
rect 430 429 756 431
rect 67 428 756 429
rect 71 422 83 423
rect 71 420 73 422
rect 75 420 83 422
rect 71 417 83 420
rect 71 415 75 417
rect 71 413 73 415
rect 71 390 75 413
rect 183 421 196 422
rect 183 419 193 421
rect 195 419 196 421
rect 183 418 196 419
rect 284 418 297 422
rect 415 422 427 423
rect 386 418 399 422
rect 95 413 117 415
rect 191 416 196 418
rect 191 414 192 416
rect 194 414 196 416
rect 95 411 114 413
rect 116 411 117 413
rect 95 409 107 411
rect 71 388 76 390
rect 71 386 73 388
rect 75 386 76 388
rect 71 381 76 386
rect 87 399 91 407
rect 87 397 99 399
rect 87 395 90 397
rect 92 396 99 397
rect 92 395 93 396
rect 87 394 93 395
rect 95 394 99 396
rect 87 393 99 394
rect 103 397 107 409
rect 105 395 107 397
rect 103 393 107 395
rect 111 406 117 411
rect 111 404 114 406
rect 116 404 117 406
rect 111 402 117 404
rect 71 379 73 381
rect 75 379 76 381
rect 71 377 76 379
rect 111 382 115 402
rect 127 405 165 406
rect 127 403 162 405
rect 164 403 165 405
rect 127 402 165 403
rect 160 399 165 402
rect 135 397 150 398
rect 135 395 139 397
rect 141 395 146 397
rect 148 395 150 397
rect 135 394 150 395
rect 160 397 168 399
rect 160 395 165 397
rect 167 395 168 397
rect 144 388 148 394
rect 160 393 168 395
rect 191 409 196 414
rect 191 407 192 409
rect 194 407 196 409
rect 191 405 196 407
rect 144 386 145 388
rect 147 386 148 388
rect 144 385 148 386
rect 111 381 133 382
rect 111 379 114 381
rect 116 379 133 381
rect 111 378 133 379
rect 192 383 196 405
rect 191 381 196 383
rect 191 379 192 381
rect 194 379 196 381
rect 191 377 196 379
rect 212 413 218 415
rect 292 416 297 418
rect 292 414 293 416
rect 295 414 297 416
rect 212 411 215 413
rect 217 411 218 413
rect 212 406 218 411
rect 212 404 215 406
rect 217 404 218 406
rect 212 402 218 404
rect 212 382 216 402
rect 228 405 266 406
rect 228 403 250 405
rect 252 403 266 405
rect 228 402 266 403
rect 261 399 266 402
rect 236 397 251 398
rect 236 395 240 397
rect 242 395 247 397
rect 249 395 251 397
rect 236 394 251 395
rect 261 397 269 399
rect 261 395 266 397
rect 268 395 269 397
rect 245 385 249 394
rect 261 393 269 395
rect 292 409 297 414
rect 292 407 293 409
rect 295 407 297 409
rect 292 405 297 407
rect 212 381 234 382
rect 212 379 215 381
rect 217 379 234 381
rect 212 378 234 379
rect 293 383 297 405
rect 292 381 297 383
rect 292 379 293 381
rect 295 379 297 381
rect 292 377 297 379
rect 314 413 320 415
rect 394 416 399 418
rect 394 414 395 416
rect 397 414 399 416
rect 314 411 317 413
rect 319 411 320 413
rect 314 406 320 411
rect 314 404 317 406
rect 319 404 320 406
rect 314 402 320 404
rect 314 382 318 402
rect 330 405 368 406
rect 330 403 331 405
rect 333 403 368 405
rect 330 402 368 403
rect 363 399 368 402
rect 338 397 353 398
rect 338 395 342 397
rect 344 395 349 397
rect 351 395 353 397
rect 338 394 353 395
rect 363 397 371 399
rect 363 395 368 397
rect 370 395 371 397
rect 347 388 351 394
rect 363 393 371 395
rect 394 409 399 414
rect 394 407 395 409
rect 397 407 399 409
rect 394 405 399 407
rect 347 386 348 388
rect 350 386 351 388
rect 347 385 351 386
rect 314 381 336 382
rect 314 379 317 381
rect 319 379 336 381
rect 314 378 336 379
rect 395 383 399 405
rect 394 381 399 383
rect 394 379 395 381
rect 397 379 399 381
rect 394 377 399 379
rect 415 420 417 422
rect 419 420 427 422
rect 415 417 427 420
rect 415 415 419 417
rect 415 413 417 415
rect 415 397 419 413
rect 539 418 552 422
rect 640 418 653 422
rect 739 418 752 422
rect 415 395 416 397
rect 418 395 419 397
rect 415 390 419 395
rect 439 413 473 415
rect 547 416 552 418
rect 547 414 548 416
rect 550 414 552 416
rect 439 411 470 413
rect 472 411 473 413
rect 439 409 451 411
rect 415 388 420 390
rect 415 386 417 388
rect 419 386 420 388
rect 415 381 420 386
rect 431 399 435 407
rect 431 397 443 399
rect 431 395 434 397
rect 436 396 443 397
rect 436 395 439 396
rect 431 394 439 395
rect 441 394 443 396
rect 431 393 443 394
rect 447 397 451 409
rect 449 395 451 397
rect 447 393 451 395
rect 467 406 473 411
rect 467 404 470 406
rect 472 404 473 406
rect 467 402 473 404
rect 415 379 417 381
rect 419 379 420 381
rect 415 377 420 379
rect 467 382 471 402
rect 483 405 521 406
rect 483 403 484 405
rect 486 403 521 405
rect 483 402 521 403
rect 516 399 521 402
rect 491 397 506 398
rect 491 395 495 397
rect 497 395 502 397
rect 504 395 506 397
rect 491 394 506 395
rect 516 397 524 399
rect 516 395 521 397
rect 523 395 524 397
rect 500 385 504 394
rect 516 393 524 395
rect 547 409 552 414
rect 547 407 548 409
rect 550 407 552 409
rect 547 405 552 407
rect 467 381 489 382
rect 467 379 470 381
rect 472 379 489 381
rect 467 378 489 379
rect 548 383 552 405
rect 547 381 552 383
rect 544 380 548 381
rect 544 378 545 380
rect 547 379 548 380
rect 550 379 552 381
rect 547 378 552 379
rect 568 413 574 415
rect 648 416 653 418
rect 648 414 649 416
rect 651 414 653 416
rect 568 411 571 413
rect 573 411 574 413
rect 568 406 574 411
rect 568 404 571 406
rect 573 404 574 406
rect 568 402 574 404
rect 568 388 572 402
rect 584 405 622 406
rect 584 403 585 405
rect 587 403 622 405
rect 584 402 622 403
rect 617 399 622 402
rect 592 397 607 398
rect 592 395 596 397
rect 598 395 603 397
rect 605 395 607 397
rect 592 394 607 395
rect 617 397 625 399
rect 617 395 622 397
rect 624 395 625 397
rect 568 386 569 388
rect 571 386 572 388
rect 568 382 572 386
rect 601 388 605 394
rect 617 393 625 395
rect 648 409 653 414
rect 648 407 649 409
rect 651 407 653 409
rect 648 405 653 407
rect 649 396 653 405
rect 649 394 650 396
rect 652 394 653 396
rect 601 386 602 388
rect 604 386 605 388
rect 601 385 605 386
rect 568 381 590 382
rect 568 379 571 381
rect 573 379 590 381
rect 568 378 590 379
rect 649 383 653 394
rect 648 381 653 383
rect 648 379 649 381
rect 651 379 653 381
rect 544 377 552 378
rect 648 377 653 379
rect 667 413 673 415
rect 747 416 752 418
rect 747 414 748 416
rect 750 414 752 416
rect 667 411 670 413
rect 672 411 673 413
rect 667 406 673 411
rect 667 404 670 406
rect 672 404 673 406
rect 667 402 673 404
rect 667 388 671 402
rect 683 405 721 406
rect 683 403 684 405
rect 686 403 721 405
rect 683 402 721 403
rect 716 399 721 402
rect 691 397 706 398
rect 691 395 692 397
rect 694 395 695 397
rect 697 395 702 397
rect 704 395 706 397
rect 691 394 706 395
rect 716 397 724 399
rect 716 395 721 397
rect 723 395 724 397
rect 667 386 668 388
rect 670 386 671 388
rect 667 382 671 386
rect 700 385 704 394
rect 716 393 724 395
rect 747 409 752 414
rect 747 407 748 409
rect 750 407 752 409
rect 747 405 752 407
rect 667 381 689 382
rect 667 379 670 381
rect 672 379 689 381
rect 667 378 689 379
rect 748 383 752 405
rect 747 381 752 383
rect 747 379 748 381
rect 750 379 752 381
rect 747 377 752 379
rect 67 371 756 372
rect 67 369 444 371
rect 446 369 756 371
rect 67 366 756 369
rect 64 365 756 366
rect 64 363 65 365
rect 67 364 193 365
rect 67 363 129 364
rect 64 362 129 363
rect 131 363 193 364
rect 195 363 257 365
rect 259 363 320 365
rect 322 363 356 365
rect 358 363 387 365
rect 389 364 606 365
rect 389 363 428 364
rect 131 362 428 363
rect 430 362 459 364
rect 461 362 516 364
rect 518 363 606 364
rect 608 363 709 365
rect 711 363 753 365
rect 755 363 756 365
rect 518 362 756 363
rect 67 359 756 362
rect 67 357 190 359
rect 192 357 444 359
rect 446 357 756 359
rect 67 356 756 357
rect 72 349 94 350
rect 72 347 75 349
rect 77 347 91 349
rect 93 347 94 349
rect 72 346 94 347
rect 152 349 157 351
rect 152 347 153 349
rect 155 347 157 349
rect 72 326 76 346
rect 105 341 109 343
rect 105 339 106 341
rect 108 339 109 341
rect 72 324 78 326
rect 72 322 75 324
rect 77 322 78 324
rect 72 317 78 322
rect 72 315 75 317
rect 77 315 78 317
rect 72 313 78 315
rect 105 334 109 339
rect 152 345 157 347
rect 96 333 111 334
rect 96 331 100 333
rect 102 331 107 333
rect 109 331 111 333
rect 96 330 111 331
rect 121 333 129 335
rect 121 331 126 333
rect 128 331 129 333
rect 121 329 129 331
rect 121 326 126 329
rect 88 325 126 326
rect 88 323 123 325
rect 125 323 126 325
rect 88 322 126 323
rect 153 323 157 345
rect 152 321 157 323
rect 152 319 153 321
rect 155 319 157 321
rect 152 314 157 319
rect 152 312 153 314
rect 155 312 157 314
rect 152 310 157 312
rect 144 306 157 310
rect 161 349 166 351
rect 161 347 163 349
rect 165 347 166 349
rect 161 342 166 347
rect 213 349 235 350
rect 213 347 216 349
rect 218 347 235 349
rect 213 346 235 347
rect 293 349 298 351
rect 293 347 294 349
rect 296 347 298 349
rect 161 340 163 342
rect 165 340 166 342
rect 161 338 166 340
rect 161 315 165 338
rect 213 335 217 346
rect 246 342 250 343
rect 246 340 247 342
rect 249 340 250 342
rect 177 334 189 335
rect 177 333 185 334
rect 177 331 180 333
rect 182 332 185 333
rect 187 332 189 334
rect 182 331 189 332
rect 177 329 189 331
rect 177 321 181 329
rect 193 333 217 335
rect 195 331 217 333
rect 193 319 197 331
rect 161 313 163 315
rect 161 311 165 313
rect 161 308 173 311
rect 161 306 163 308
rect 165 306 173 308
rect 161 305 173 306
rect 185 313 197 319
rect 213 326 217 331
rect 213 324 219 326
rect 213 322 216 324
rect 218 322 219 324
rect 213 317 219 322
rect 213 315 216 317
rect 218 315 219 317
rect 213 313 219 315
rect 246 334 250 340
rect 293 345 298 347
rect 294 341 298 345
rect 294 339 295 341
rect 297 339 298 341
rect 237 333 252 334
rect 237 331 241 333
rect 243 331 248 333
rect 250 331 252 333
rect 237 330 252 331
rect 262 333 270 335
rect 262 331 267 333
rect 269 331 270 333
rect 262 329 270 331
rect 262 326 267 329
rect 229 322 267 326
rect 294 323 298 339
rect 293 321 298 323
rect 293 319 294 321
rect 296 319 298 321
rect 293 314 298 319
rect 293 312 294 314
rect 296 312 298 314
rect 293 310 298 312
rect 285 306 298 310
rect 314 349 319 351
rect 314 347 316 349
rect 318 347 319 349
rect 314 345 319 347
rect 314 323 318 345
rect 377 349 399 350
rect 377 347 378 349
rect 380 347 394 349
rect 396 347 399 349
rect 377 346 399 347
rect 362 341 366 343
rect 362 339 363 341
rect 365 339 366 341
rect 314 321 319 323
rect 314 319 316 321
rect 318 319 319 321
rect 314 314 319 319
rect 342 333 350 335
rect 362 334 366 339
rect 342 331 343 333
rect 345 331 350 333
rect 342 329 350 331
rect 360 333 375 334
rect 360 331 362 333
rect 364 331 369 333
rect 371 331 375 333
rect 360 330 375 331
rect 345 326 350 329
rect 345 325 383 326
rect 345 323 380 325
rect 382 323 383 325
rect 345 322 383 323
rect 395 326 399 346
rect 393 324 399 326
rect 393 322 394 324
rect 396 322 399 324
rect 393 317 399 322
rect 393 315 394 317
rect 396 315 399 317
rect 314 312 316 314
rect 318 312 319 314
rect 314 310 319 312
rect 393 313 399 315
rect 415 349 420 351
rect 415 347 417 349
rect 419 347 420 349
rect 415 342 420 347
rect 467 349 489 350
rect 467 347 470 349
rect 472 347 489 349
rect 467 346 489 347
rect 547 349 552 351
rect 547 347 548 349
rect 550 347 552 349
rect 415 340 417 342
rect 419 340 420 342
rect 415 338 420 340
rect 415 325 419 338
rect 415 323 416 325
rect 418 323 419 325
rect 415 315 419 323
rect 431 334 443 335
rect 431 333 439 334
rect 431 331 434 333
rect 436 332 439 333
rect 441 332 443 334
rect 436 331 443 332
rect 431 329 443 331
rect 431 321 435 329
rect 447 333 451 335
rect 449 331 451 333
rect 447 319 451 331
rect 415 313 417 315
rect 415 311 419 313
rect 314 309 327 310
rect 314 307 324 309
rect 326 307 327 309
rect 314 306 327 307
rect 415 308 427 311
rect 415 306 417 308
rect 419 306 427 308
rect 415 305 427 306
rect 439 317 451 319
rect 467 326 471 346
rect 467 324 473 326
rect 467 322 470 324
rect 472 322 473 324
rect 467 317 473 322
rect 439 315 470 317
rect 472 315 473 317
rect 439 313 473 315
rect 500 334 504 343
rect 547 345 552 347
rect 491 333 506 334
rect 491 331 495 333
rect 497 331 502 333
rect 504 331 506 333
rect 491 330 506 331
rect 516 333 524 335
rect 516 331 521 333
rect 523 331 524 333
rect 516 329 524 331
rect 516 326 521 329
rect 483 325 521 326
rect 483 323 518 325
rect 520 323 521 325
rect 483 322 521 323
rect 548 323 552 345
rect 547 321 552 323
rect 547 319 548 321
rect 550 319 552 321
rect 547 314 552 319
rect 547 312 548 314
rect 550 312 552 314
rect 568 349 590 350
rect 568 347 571 349
rect 573 347 590 349
rect 568 346 590 347
rect 648 349 653 351
rect 648 347 649 349
rect 651 347 653 349
rect 568 342 572 346
rect 568 340 569 342
rect 571 340 572 342
rect 568 326 572 340
rect 601 342 605 343
rect 601 340 602 342
rect 604 340 605 342
rect 568 324 574 326
rect 568 322 571 324
rect 573 322 574 324
rect 568 317 574 322
rect 568 315 571 317
rect 573 315 574 317
rect 568 313 574 315
rect 601 334 605 340
rect 648 345 653 347
rect 592 333 607 334
rect 592 331 596 333
rect 598 331 603 333
rect 605 331 607 333
rect 592 330 607 331
rect 617 333 625 335
rect 617 331 622 333
rect 624 331 625 333
rect 617 329 625 331
rect 617 326 622 329
rect 649 334 653 345
rect 649 332 650 334
rect 652 332 653 334
rect 584 324 619 326
rect 621 324 622 326
rect 584 322 622 324
rect 649 323 653 332
rect 648 321 653 323
rect 648 319 649 321
rect 651 319 653 321
rect 648 314 653 319
rect 547 310 552 312
rect 648 312 649 314
rect 651 312 653 314
rect 667 349 689 350
rect 667 347 670 349
rect 672 347 689 349
rect 667 346 689 347
rect 747 349 752 351
rect 747 347 748 349
rect 750 347 752 349
rect 667 342 671 346
rect 667 340 668 342
rect 670 340 671 342
rect 667 326 671 340
rect 700 342 704 343
rect 700 340 701 342
rect 703 340 704 342
rect 667 324 673 326
rect 667 322 670 324
rect 672 322 673 324
rect 667 317 673 322
rect 667 315 670 317
rect 672 315 673 317
rect 667 313 673 315
rect 700 334 704 340
rect 747 345 752 347
rect 691 333 706 334
rect 691 331 695 333
rect 697 331 702 333
rect 704 331 706 333
rect 691 330 706 331
rect 716 333 724 335
rect 716 331 721 333
rect 723 331 724 333
rect 716 329 724 331
rect 716 326 721 329
rect 683 325 721 326
rect 683 323 718 325
rect 720 323 721 325
rect 683 322 721 323
rect 748 323 752 345
rect 747 321 752 323
rect 747 319 748 321
rect 750 319 752 321
rect 747 314 752 319
rect 648 310 653 312
rect 747 312 748 314
rect 750 312 752 314
rect 747 310 752 312
rect 539 306 552 310
rect 640 306 653 310
rect 739 306 752 310
rect 67 299 755 300
rect 67 297 174 299
rect 176 297 428 299
rect 430 297 755 299
rect 67 294 755 297
rect 64 293 109 294
rect 64 291 65 293
rect 67 292 109 293
rect 111 293 755 294
rect 111 292 146 293
rect 67 291 146 292
rect 148 291 217 293
rect 219 291 282 293
rect 284 291 335 293
rect 337 292 403 293
rect 337 291 370 292
rect 64 290 370 291
rect 372 291 403 292
rect 405 291 449 293
rect 451 291 494 293
rect 496 292 752 293
rect 496 291 567 292
rect 372 290 567 291
rect 569 290 632 292
rect 634 291 752 292
rect 754 291 755 293
rect 634 290 755 291
rect 67 287 755 290
rect 67 285 84 287
rect 86 285 427 287
rect 429 285 755 287
rect 67 284 755 285
rect 71 278 83 279
rect 71 276 73 278
rect 75 276 83 278
rect 71 273 83 276
rect 71 271 75 273
rect 71 269 73 271
rect 71 246 75 269
rect 183 274 196 278
rect 284 274 297 278
rect 414 278 426 279
rect 385 274 398 278
rect 95 269 117 271
rect 191 272 196 274
rect 191 270 192 272
rect 194 270 196 272
rect 95 267 114 269
rect 116 267 117 269
rect 95 265 107 267
rect 71 244 76 246
rect 71 242 73 244
rect 75 242 76 244
rect 71 237 76 242
rect 87 255 91 263
rect 87 253 99 255
rect 87 251 90 253
rect 92 252 99 253
rect 92 251 95 252
rect 87 250 95 251
rect 97 250 99 252
rect 87 249 99 250
rect 103 253 107 265
rect 105 251 107 253
rect 103 249 107 251
rect 111 262 117 267
rect 111 260 114 262
rect 116 260 117 262
rect 111 258 117 260
rect 71 235 73 237
rect 75 235 76 237
rect 71 233 76 235
rect 111 238 115 258
rect 127 261 165 262
rect 127 259 128 261
rect 130 259 165 261
rect 127 258 165 259
rect 160 255 165 258
rect 135 253 150 254
rect 135 251 139 253
rect 141 251 146 253
rect 148 251 150 253
rect 135 250 150 251
rect 160 253 168 255
rect 160 251 165 253
rect 167 251 168 253
rect 144 241 148 250
rect 160 249 168 251
rect 191 265 196 270
rect 191 263 192 265
rect 194 263 196 265
rect 191 261 196 263
rect 111 237 133 238
rect 111 235 114 237
rect 116 235 133 237
rect 111 234 133 235
rect 192 239 196 261
rect 191 237 196 239
rect 191 235 192 237
rect 194 235 196 237
rect 191 233 196 235
rect 212 269 218 271
rect 292 272 297 274
rect 292 270 293 272
rect 295 270 297 272
rect 212 267 215 269
rect 217 267 218 269
rect 212 262 218 267
rect 212 260 215 262
rect 217 260 218 262
rect 212 258 218 260
rect 212 244 216 258
rect 228 261 266 262
rect 228 259 229 261
rect 231 259 266 261
rect 228 258 266 259
rect 261 255 266 258
rect 236 253 251 254
rect 236 251 240 253
rect 242 251 247 253
rect 249 251 251 253
rect 236 250 251 251
rect 261 253 269 255
rect 261 251 266 253
rect 268 251 269 253
rect 212 242 213 244
rect 215 242 216 244
rect 212 238 216 242
rect 245 244 249 250
rect 261 249 269 251
rect 292 265 297 270
rect 292 263 293 265
rect 295 263 297 265
rect 292 261 297 263
rect 293 252 297 261
rect 293 250 294 252
rect 296 250 297 252
rect 245 242 246 244
rect 248 242 249 244
rect 245 241 249 242
rect 212 237 234 238
rect 212 235 215 237
rect 217 235 234 237
rect 212 234 234 235
rect 293 239 297 250
rect 292 237 297 239
rect 292 235 293 237
rect 295 235 297 237
rect 292 233 297 235
rect 313 269 319 271
rect 393 272 398 274
rect 393 270 394 272
rect 396 270 398 272
rect 313 267 316 269
rect 318 267 319 269
rect 313 262 319 267
rect 313 260 316 262
rect 318 260 319 262
rect 313 258 319 260
rect 313 244 317 258
rect 329 261 367 262
rect 329 259 330 261
rect 332 259 367 261
rect 329 258 367 259
rect 362 255 367 258
rect 337 253 352 254
rect 337 251 341 253
rect 343 251 348 253
rect 350 251 352 253
rect 337 250 352 251
rect 362 253 370 255
rect 362 251 367 253
rect 369 251 370 253
rect 346 249 350 250
rect 362 249 370 251
rect 313 242 314 244
rect 316 242 317 244
rect 346 247 347 249
rect 349 247 350 249
rect 313 238 317 242
rect 346 241 350 247
rect 393 265 398 270
rect 393 263 394 265
rect 396 263 398 265
rect 393 261 398 263
rect 313 237 335 238
rect 313 235 316 237
rect 318 235 335 237
rect 313 234 335 235
rect 394 239 398 261
rect 393 237 398 239
rect 393 235 394 237
rect 396 235 398 237
rect 393 233 398 235
rect 414 276 416 278
rect 418 276 426 278
rect 414 273 426 276
rect 414 271 418 273
rect 414 269 416 271
rect 414 249 418 269
rect 538 274 551 278
rect 639 274 652 278
rect 738 274 751 278
rect 414 247 415 249
rect 417 247 418 249
rect 414 246 418 247
rect 438 269 472 271
rect 546 272 551 274
rect 546 270 547 272
rect 549 270 551 272
rect 438 267 469 269
rect 471 267 472 269
rect 438 265 450 267
rect 414 244 419 246
rect 414 242 416 244
rect 418 242 419 244
rect 414 237 419 242
rect 430 255 434 263
rect 430 253 442 255
rect 430 251 433 253
rect 435 252 442 253
rect 435 251 438 252
rect 430 250 438 251
rect 440 250 442 252
rect 430 249 442 250
rect 446 253 450 265
rect 448 251 450 253
rect 446 249 450 251
rect 466 262 472 267
rect 466 260 469 262
rect 471 260 472 262
rect 466 258 472 260
rect 414 235 416 237
rect 418 235 419 237
rect 414 233 419 235
rect 466 238 470 258
rect 482 261 520 262
rect 482 259 483 261
rect 485 259 520 261
rect 482 258 520 259
rect 515 255 520 258
rect 490 253 505 254
rect 490 251 494 253
rect 496 251 501 253
rect 503 251 505 253
rect 490 250 505 251
rect 515 253 523 255
rect 515 251 520 253
rect 522 251 523 253
rect 499 241 503 250
rect 515 249 523 251
rect 546 265 551 270
rect 546 263 547 265
rect 549 263 551 265
rect 546 261 551 263
rect 466 237 488 238
rect 466 235 469 237
rect 471 235 488 237
rect 466 234 488 235
rect 547 239 551 261
rect 546 237 551 239
rect 546 235 547 237
rect 549 235 551 237
rect 546 233 551 235
rect 567 269 573 271
rect 647 272 652 274
rect 647 270 648 272
rect 650 270 652 272
rect 567 267 570 269
rect 572 267 573 269
rect 567 262 573 267
rect 567 260 570 262
rect 572 260 573 262
rect 567 258 573 260
rect 567 244 571 258
rect 583 261 621 262
rect 583 259 584 261
rect 586 259 621 261
rect 583 258 621 259
rect 616 255 621 258
rect 591 253 606 254
rect 591 251 595 253
rect 597 251 602 253
rect 604 251 606 253
rect 591 250 606 251
rect 616 253 624 255
rect 616 251 621 253
rect 623 251 624 253
rect 567 242 568 244
rect 570 242 571 244
rect 567 238 571 242
rect 600 244 604 250
rect 616 249 624 251
rect 647 265 652 270
rect 647 263 648 265
rect 650 263 652 265
rect 647 261 652 263
rect 648 252 652 261
rect 648 250 649 252
rect 651 250 652 252
rect 600 242 601 244
rect 603 242 604 244
rect 600 241 604 242
rect 567 237 589 238
rect 567 235 570 237
rect 572 235 589 237
rect 567 234 589 235
rect 648 239 652 250
rect 647 237 652 239
rect 647 235 648 237
rect 650 235 652 237
rect 647 233 652 235
rect 666 269 672 271
rect 746 272 751 274
rect 746 270 747 272
rect 749 270 751 272
rect 666 267 669 269
rect 671 267 672 269
rect 666 262 672 267
rect 666 260 669 262
rect 671 260 672 262
rect 666 258 672 260
rect 666 244 670 258
rect 682 261 720 262
rect 682 259 683 261
rect 685 259 720 261
rect 682 258 720 259
rect 715 255 720 258
rect 690 253 705 254
rect 690 251 691 253
rect 693 251 694 253
rect 696 251 701 253
rect 703 251 705 253
rect 690 250 705 251
rect 715 253 723 255
rect 715 251 720 253
rect 722 251 723 253
rect 666 242 667 244
rect 669 242 670 244
rect 666 238 670 242
rect 699 241 703 250
rect 715 249 723 251
rect 746 265 751 270
rect 746 263 747 265
rect 749 263 751 265
rect 746 261 751 263
rect 666 237 688 238
rect 666 235 669 237
rect 671 235 688 237
rect 666 234 688 235
rect 747 239 751 261
rect 746 237 751 239
rect 746 235 747 237
rect 749 235 751 237
rect 746 233 751 235
rect 67 227 755 228
rect 67 225 100 227
rect 102 225 443 227
rect 445 225 755 227
rect 67 223 68 225
rect 70 223 709 225
rect 711 223 752 225
rect 754 223 755 225
rect 67 220 755 223
rect 128 218 129 220
rect 131 218 132 220
rect 128 217 132 218
rect 192 218 193 220
rect 195 218 196 220
rect 192 217 196 218
rect 256 218 257 220
rect 259 218 260 220
rect 256 217 260 218
rect 319 218 320 220
rect 322 218 323 220
rect 319 217 323 218
rect 355 218 356 220
rect 358 218 359 220
rect 355 217 359 218
rect 386 218 387 220
rect 389 218 390 220
rect 386 217 390 218
rect 427 218 428 220
rect 430 218 431 220
rect 427 217 431 218
rect 458 218 459 220
rect 461 218 462 220
rect 458 217 462 218
rect 515 218 516 220
rect 518 218 519 220
rect 515 217 519 218
rect 605 218 606 220
rect 608 218 609 220
rect 605 217 609 218
<< alu2 >>
rect 402 581 406 582
rect 402 579 403 581
rect 405 579 406 581
rect 107 578 111 579
rect 402 578 406 579
rect 448 581 452 582
rect 448 579 449 581
rect 451 579 452 581
rect 448 578 452 579
rect 493 581 497 582
rect 493 579 494 581
rect 496 579 497 581
rect 493 578 497 579
rect 566 581 570 582
rect 566 579 567 581
rect 569 579 570 581
rect 566 578 570 579
rect 752 578 756 579
rect 67 577 71 578
rect 67 575 68 577
rect 70 575 71 577
rect 107 576 108 578
rect 110 576 111 578
rect 107 575 111 576
rect 145 577 149 578
rect 145 575 146 577
rect 148 575 149 577
rect 67 574 71 575
rect 145 574 149 575
rect 216 577 220 578
rect 216 575 217 577
rect 219 575 220 577
rect 216 574 220 575
rect 281 577 285 578
rect 281 575 282 577
rect 284 575 285 577
rect 281 574 285 575
rect 334 577 338 578
rect 334 575 335 577
rect 337 575 338 577
rect 334 574 338 575
rect 369 577 373 578
rect 369 575 370 577
rect 372 575 373 577
rect 369 574 373 575
rect 631 577 635 578
rect 631 575 632 577
rect 634 575 635 577
rect 752 576 753 578
rect 755 576 756 578
rect 752 575 756 576
rect 631 574 635 575
rect 400 573 600 574
rect 400 571 401 573
rect 403 571 597 573
rect 599 571 600 573
rect 400 570 600 571
rect 102 565 171 566
rect 102 563 103 565
rect 105 563 168 565
rect 170 563 171 565
rect 102 562 171 563
rect 313 565 382 566
rect 313 563 314 565
rect 316 563 379 565
rect 381 563 382 565
rect 313 562 382 563
rect 483 565 552 566
rect 483 563 484 565
rect 486 563 549 565
rect 551 563 552 565
rect 483 562 552 563
rect 618 565 687 566
rect 618 563 619 565
rect 621 563 684 565
rect 686 563 687 565
rect 618 562 687 563
rect 111 557 543 558
rect 111 555 112 557
rect 114 555 540 557
rect 542 555 543 557
rect 111 554 543 555
rect 80 549 115 550
rect 80 547 81 549
rect 83 547 112 549
rect 114 547 115 549
rect 80 546 115 547
rect 167 549 171 550
rect 167 547 168 549
rect 170 547 171 549
rect 167 546 171 547
rect 313 549 317 550
rect 313 547 314 549
rect 316 547 317 549
rect 313 546 317 547
rect 369 549 404 550
rect 369 547 370 549
rect 372 547 401 549
rect 403 547 404 549
rect 369 546 404 547
rect 483 549 487 550
rect 483 547 484 549
rect 486 547 487 549
rect 483 546 487 547
rect 539 549 574 550
rect 539 547 540 549
rect 542 547 571 549
rect 573 547 574 549
rect 539 546 574 547
rect 596 549 631 550
rect 596 547 597 549
rect 599 547 628 549
rect 630 547 631 549
rect 596 546 631 547
rect 683 549 687 550
rect 683 547 684 549
rect 686 547 687 549
rect 683 546 687 547
rect 78 541 406 542
rect 78 539 79 541
rect 81 539 403 541
rect 405 539 406 541
rect 78 538 406 539
rect 532 540 638 541
rect 532 538 533 540
rect 535 538 635 540
rect 637 538 638 540
rect 532 537 638 538
rect 78 532 82 533
rect 78 530 79 532
rect 81 530 82 532
rect 78 529 82 530
rect 118 532 122 533
rect 118 530 119 532
rect 121 530 122 532
rect 118 529 122 530
rect 184 532 188 533
rect 184 530 185 532
rect 187 530 188 532
rect 184 529 188 530
rect 296 532 300 533
rect 296 530 297 532
rect 299 530 300 532
rect 296 529 300 530
rect 362 532 366 533
rect 362 530 363 532
rect 365 530 366 532
rect 362 529 366 530
rect 402 532 406 533
rect 402 530 403 532
rect 405 530 406 532
rect 402 529 406 530
rect 466 532 470 533
rect 466 530 467 532
rect 469 530 470 532
rect 466 529 470 530
rect 532 532 536 533
rect 532 530 533 532
rect 535 530 536 532
rect 532 529 536 530
rect 572 532 576 533
rect 572 530 573 532
rect 575 530 576 532
rect 572 529 576 530
rect 594 532 598 533
rect 594 530 595 532
rect 597 530 598 532
rect 594 529 598 530
rect 634 532 638 533
rect 634 530 635 532
rect 637 530 638 532
rect 634 529 638 530
rect 700 532 704 533
rect 700 530 701 532
rect 703 530 704 532
rect 700 529 704 530
rect 169 525 173 526
rect 142 524 150 525
rect 142 522 143 524
rect 145 522 147 524
rect 149 522 150 524
rect 169 523 170 525
rect 172 523 173 525
rect 169 522 173 523
rect 231 525 240 526
rect 231 523 232 525
rect 234 523 237 525
rect 239 523 240 525
rect 231 522 240 523
rect 249 525 253 526
rect 249 523 250 525
rect 252 523 253 525
rect 249 522 253 523
rect 311 525 315 526
rect 419 525 423 526
rect 311 523 312 525
rect 314 523 315 525
rect 311 522 315 523
rect 334 524 342 525
rect 334 522 335 524
rect 337 522 339 524
rect 341 522 342 524
rect 419 523 420 525
rect 422 523 423 525
rect 419 522 423 523
rect 481 525 485 526
rect 685 525 689 526
rect 481 523 482 525
rect 484 523 485 525
rect 481 522 485 523
rect 504 524 512 525
rect 504 522 505 524
rect 507 522 509 524
rect 511 522 512 524
rect 142 521 150 522
rect 334 521 342 522
rect 504 521 512 522
rect 658 524 666 525
rect 658 522 659 524
rect 661 522 663 524
rect 665 522 666 524
rect 685 523 686 525
rect 688 523 689 525
rect 685 522 689 523
rect 658 521 666 522
rect 67 509 71 510
rect 67 507 68 509
rect 70 507 71 509
rect 67 506 71 507
rect 128 509 132 510
rect 128 507 129 509
rect 131 507 132 509
rect 128 506 132 507
rect 192 509 196 510
rect 192 507 193 509
rect 195 507 196 509
rect 192 506 196 507
rect 256 509 260 510
rect 256 507 257 509
rect 259 507 260 509
rect 256 506 260 507
rect 319 509 323 510
rect 319 507 320 509
rect 322 507 323 509
rect 319 506 323 507
rect 354 509 358 510
rect 354 507 355 509
rect 357 507 358 509
rect 354 506 358 507
rect 386 509 390 510
rect 386 507 387 509
rect 389 507 390 509
rect 386 506 390 507
rect 427 509 431 510
rect 427 507 428 509
rect 430 507 431 509
rect 427 506 431 507
rect 458 509 462 510
rect 458 507 459 509
rect 461 507 462 509
rect 458 506 462 507
rect 515 509 519 510
rect 515 507 516 509
rect 518 507 519 509
rect 515 506 519 507
rect 605 509 609 510
rect 605 507 606 509
rect 608 507 609 509
rect 605 506 609 507
rect 708 509 712 510
rect 708 507 709 509
rect 711 507 712 509
rect 708 506 712 507
rect 752 509 756 510
rect 752 507 753 509
rect 755 507 756 509
rect 752 506 756 507
rect 142 494 188 495
rect 142 492 143 494
rect 145 492 185 494
rect 187 492 188 494
rect 142 491 188 492
rect 296 494 342 495
rect 296 492 297 494
rect 299 492 339 494
rect 341 492 342 494
rect 296 491 342 492
rect 466 494 512 495
rect 466 492 467 494
rect 469 492 509 494
rect 511 492 512 494
rect 466 491 512 492
rect 658 494 704 495
rect 658 492 659 494
rect 661 492 701 494
rect 703 492 704 494
rect 658 491 704 492
rect 78 486 82 487
rect 78 484 79 486
rect 81 484 82 486
rect 78 483 82 484
rect 118 486 366 487
rect 118 484 119 486
rect 121 484 363 486
rect 365 484 366 486
rect 118 483 366 484
rect 402 486 406 487
rect 532 486 536 487
rect 402 484 403 486
rect 405 484 406 486
rect 402 483 406 484
rect 458 485 503 486
rect 458 483 459 485
rect 461 483 500 485
rect 502 483 503 485
rect 532 484 533 486
rect 535 484 536 486
rect 532 483 536 484
rect 572 486 598 487
rect 572 484 573 486
rect 575 484 595 486
rect 597 484 598 486
rect 572 483 598 484
rect 634 486 638 487
rect 634 484 635 486
rect 637 484 638 486
rect 634 483 638 484
rect 458 482 503 483
rect 99 477 107 478
rect 99 475 100 477
rect 102 475 104 477
rect 106 475 107 477
rect 99 474 107 475
rect 169 477 179 478
rect 169 475 170 477
rect 172 475 176 477
rect 178 475 179 477
rect 169 474 179 475
rect 248 477 301 478
rect 248 475 249 477
rect 251 475 298 477
rect 300 475 301 477
rect 248 474 301 475
rect 305 477 315 478
rect 305 475 306 477
rect 308 475 312 477
rect 314 475 315 477
rect 305 474 315 475
rect 475 477 485 478
rect 475 475 476 477
rect 478 475 482 477
rect 484 475 485 477
rect 475 474 485 475
rect 547 477 562 478
rect 547 475 548 477
rect 550 475 559 477
rect 561 475 562 477
rect 547 474 562 475
rect 685 477 695 478
rect 685 475 686 477
rect 688 475 692 477
rect 694 475 695 477
rect 685 474 695 475
rect 80 469 115 470
rect 80 467 81 469
rect 83 467 108 469
rect 110 467 112 469
rect 114 467 115 469
rect 80 466 115 467
rect 146 469 171 470
rect 146 467 147 469
rect 149 467 168 469
rect 170 467 171 469
rect 146 466 171 467
rect 208 469 262 470
rect 208 467 209 469
rect 211 467 259 469
rect 261 467 262 469
rect 208 466 262 467
rect 313 469 338 470
rect 313 467 314 469
rect 316 467 335 469
rect 337 467 338 469
rect 313 466 338 467
rect 369 469 404 470
rect 369 467 370 469
rect 372 467 401 469
rect 403 467 404 469
rect 369 466 404 467
rect 483 469 508 470
rect 483 467 484 469
rect 486 467 505 469
rect 507 467 508 469
rect 483 466 508 467
rect 539 469 574 470
rect 539 467 540 469
rect 542 467 571 469
rect 573 467 574 469
rect 539 466 574 467
rect 596 469 631 470
rect 596 467 597 469
rect 599 467 628 469
rect 630 467 631 469
rect 596 466 631 467
rect 662 469 687 470
rect 662 467 663 469
rect 665 467 684 469
rect 686 467 687 469
rect 662 466 687 467
rect 409 465 423 466
rect 409 463 410 465
rect 412 463 420 465
rect 422 463 423 465
rect 409 462 423 463
rect 153 461 157 462
rect 153 459 154 461
rect 156 459 157 461
rect 258 461 331 462
rect 258 459 259 461
rect 261 459 328 461
rect 330 459 331 461
rect 153 458 157 459
rect 227 458 235 459
rect 227 456 228 458
rect 230 456 232 458
rect 234 456 235 458
rect 227 455 235 456
rect 249 458 253 459
rect 258 458 331 459
rect 653 461 673 462
rect 653 459 654 461
rect 656 459 670 461
rect 672 459 673 461
rect 653 458 673 459
rect 249 456 250 458
rect 252 456 253 458
rect 249 455 253 456
rect 378 456 382 457
rect 378 454 379 456
rect 381 454 382 456
rect 378 453 382 454
rect 400 456 600 457
rect 400 454 401 456
rect 403 454 597 456
rect 599 454 600 456
rect 400 453 600 454
rect 739 453 743 454
rect 739 451 740 453
rect 742 451 743 453
rect 739 450 743 451
rect 107 448 543 449
rect 107 446 108 448
rect 110 446 540 448
rect 542 446 543 448
rect 107 445 543 446
rect 752 438 756 439
rect 107 437 111 438
rect 67 436 71 437
rect 67 434 68 436
rect 70 434 71 436
rect 107 435 108 437
rect 110 435 111 437
rect 107 434 111 435
rect 145 437 149 438
rect 145 435 146 437
rect 148 435 149 437
rect 145 434 149 435
rect 216 437 220 438
rect 216 435 217 437
rect 219 435 220 437
rect 216 434 220 435
rect 281 437 285 438
rect 281 435 282 437
rect 284 435 285 437
rect 281 434 285 435
rect 334 437 338 438
rect 448 437 452 438
rect 334 435 335 437
rect 337 435 338 437
rect 334 434 338 435
rect 369 436 373 437
rect 369 434 370 436
rect 372 434 373 436
rect 67 433 71 434
rect 369 433 373 434
rect 401 436 405 437
rect 401 434 402 436
rect 404 434 405 436
rect 448 435 449 437
rect 451 435 452 437
rect 448 434 452 435
rect 493 437 497 438
rect 493 435 494 437
rect 496 435 497 437
rect 493 434 497 435
rect 566 436 570 437
rect 566 434 567 436
rect 569 434 570 436
rect 401 433 405 434
rect 566 433 570 434
rect 631 436 635 437
rect 631 434 632 436
rect 634 434 635 436
rect 752 436 753 438
rect 755 436 756 438
rect 752 435 756 436
rect 631 433 635 434
rect 192 421 334 422
rect 192 419 193 421
rect 195 419 331 421
rect 333 419 334 421
rect 192 418 334 419
rect 378 421 687 422
rect 378 419 379 421
rect 381 419 684 421
rect 686 419 687 421
rect 378 418 687 419
rect 297 413 487 414
rect 297 411 298 413
rect 300 411 484 413
rect 486 411 487 413
rect 297 410 487 411
rect 558 413 695 414
rect 558 411 559 413
rect 561 411 692 413
rect 694 411 695 413
rect 558 410 695 411
rect 161 405 204 406
rect 161 403 162 405
rect 164 403 201 405
rect 203 403 204 405
rect 161 402 204 403
rect 249 405 253 406
rect 249 403 250 405
rect 252 403 253 405
rect 249 402 253 403
rect 330 405 334 406
rect 330 403 331 405
rect 333 403 334 405
rect 330 402 334 403
rect 358 405 462 406
rect 358 403 359 405
rect 361 403 459 405
rect 461 403 462 405
rect 358 402 462 403
rect 483 405 487 406
rect 483 403 484 405
rect 486 403 487 405
rect 483 402 487 403
rect 584 405 588 406
rect 584 403 585 405
rect 587 403 588 405
rect 584 402 588 403
rect 683 405 687 406
rect 683 403 684 405
rect 686 403 687 405
rect 683 402 687 403
rect 246 397 419 398
rect 501 397 505 398
rect 691 397 695 398
rect 92 396 96 397
rect 92 394 93 396
rect 95 394 96 396
rect 92 393 96 394
rect 153 396 165 397
rect 153 394 154 396
rect 156 394 162 396
rect 164 394 165 396
rect 246 395 247 397
rect 249 395 416 397
rect 418 395 419 397
rect 246 394 419 395
rect 438 396 442 397
rect 438 394 439 396
rect 441 394 442 396
rect 153 393 165 394
rect 200 389 308 390
rect 438 389 442 394
rect 501 395 502 397
rect 504 396 653 397
rect 504 395 650 396
rect 501 394 650 395
rect 652 394 653 396
rect 691 395 692 397
rect 694 395 695 397
rect 691 394 695 395
rect 501 393 653 394
rect 144 388 156 389
rect 144 386 145 388
rect 147 386 153 388
rect 155 386 156 388
rect 200 387 201 389
rect 203 387 305 389
rect 307 387 308 389
rect 200 386 308 387
rect 347 388 351 389
rect 347 386 348 388
rect 350 386 351 388
rect 144 385 156 386
rect 347 385 351 386
rect 438 388 572 389
rect 438 386 569 388
rect 571 386 572 388
rect 438 385 572 386
rect 601 388 671 389
rect 601 386 602 388
rect 604 386 668 388
rect 670 386 671 388
rect 601 385 671 386
rect 72 381 76 382
rect 72 379 73 381
rect 75 379 76 381
rect 72 378 76 379
rect 184 381 218 382
rect 184 379 185 381
rect 187 379 215 381
rect 217 379 218 381
rect 184 378 218 379
rect 245 381 296 382
rect 394 381 398 382
rect 700 381 751 382
rect 245 379 247 381
rect 249 379 293 381
rect 295 379 296 381
rect 245 378 296 379
rect 304 380 362 381
rect 304 378 305 380
rect 307 378 359 380
rect 361 378 362 380
rect 394 379 395 381
rect 397 379 398 381
rect 394 378 398 379
rect 544 380 548 381
rect 544 378 545 380
rect 547 378 548 380
rect 700 379 701 381
rect 703 379 748 381
rect 750 379 751 381
rect 700 378 751 379
rect 304 377 362 378
rect 544 377 548 378
rect 419 372 588 373
rect 419 370 420 372
rect 422 370 585 372
rect 587 370 588 372
rect 419 369 588 370
rect 64 365 68 366
rect 192 365 196 366
rect 64 363 65 365
rect 67 363 68 365
rect 64 362 68 363
rect 128 364 132 365
rect 128 362 129 364
rect 131 362 132 364
rect 192 363 193 365
rect 195 363 196 365
rect 192 362 196 363
rect 256 365 260 366
rect 256 363 257 365
rect 259 363 260 365
rect 256 362 260 363
rect 319 365 323 366
rect 319 363 320 365
rect 322 363 323 365
rect 319 362 323 363
rect 355 365 359 366
rect 355 363 356 365
rect 358 363 359 365
rect 355 362 359 363
rect 386 365 390 366
rect 605 365 609 366
rect 386 363 387 365
rect 389 363 390 365
rect 386 362 390 363
rect 427 364 431 365
rect 427 362 428 364
rect 430 362 431 364
rect 128 361 132 362
rect 427 361 431 362
rect 458 364 462 365
rect 458 362 459 364
rect 461 362 462 364
rect 458 361 462 362
rect 515 364 519 365
rect 515 362 516 364
rect 518 362 519 364
rect 605 363 606 365
rect 608 363 609 365
rect 605 362 609 363
rect 708 365 712 366
rect 708 363 709 365
rect 711 363 712 365
rect 708 362 712 363
rect 752 365 756 366
rect 752 363 753 365
rect 755 363 756 365
rect 752 362 756 363
rect 515 361 519 362
rect 90 349 94 350
rect 90 347 91 349
rect 93 347 94 349
rect 90 346 94 347
rect 152 349 156 350
rect 152 347 153 349
rect 155 347 156 349
rect 152 346 156 347
rect 347 349 381 350
rect 347 347 348 349
rect 350 347 378 349
rect 380 347 381 349
rect 347 346 381 347
rect 162 342 166 343
rect 105 341 163 342
rect 105 339 106 341
rect 108 340 163 341
rect 165 340 166 342
rect 108 339 166 340
rect 246 342 250 343
rect 438 342 572 343
rect 246 340 247 342
rect 249 340 250 342
rect 246 339 250 340
rect 294 341 366 342
rect 294 339 295 341
rect 297 339 363 341
rect 365 339 366 341
rect 105 338 166 339
rect 294 338 366 339
rect 438 340 569 342
rect 571 340 572 342
rect 438 339 572 340
rect 601 342 671 343
rect 601 340 602 342
rect 604 340 668 342
rect 670 340 671 342
rect 601 339 671 340
rect 700 342 704 343
rect 700 340 701 342
rect 703 340 704 342
rect 700 339 704 340
rect 184 334 188 335
rect 438 334 442 339
rect 184 332 185 334
rect 187 332 188 334
rect 184 331 188 332
rect 266 333 413 334
rect 266 331 267 333
rect 269 331 410 333
rect 412 331 413 333
rect 438 332 439 334
rect 441 332 442 334
rect 438 331 442 332
rect 501 334 653 335
rect 501 333 650 334
rect 501 331 502 333
rect 504 332 650 333
rect 652 332 653 334
rect 504 331 653 332
rect 266 330 413 331
rect 501 330 505 331
rect 618 326 657 327
rect 122 325 212 326
rect 122 323 123 325
rect 125 323 209 325
rect 211 323 212 325
rect 122 322 212 323
rect 379 325 419 326
rect 379 323 380 325
rect 382 323 416 325
rect 418 323 419 325
rect 379 322 419 323
rect 517 325 548 326
rect 517 323 518 325
rect 520 323 545 325
rect 547 323 548 325
rect 618 324 619 326
rect 621 324 654 326
rect 656 324 657 326
rect 618 323 657 324
rect 717 325 743 326
rect 717 323 718 325
rect 720 323 740 325
rect 742 323 743 325
rect 517 322 548 323
rect 717 322 743 323
rect 323 309 327 310
rect 323 307 324 309
rect 326 307 327 309
rect 323 306 327 307
rect 323 301 694 302
rect 323 299 324 301
rect 326 299 691 301
rect 693 299 694 301
rect 323 298 694 299
rect 108 294 112 295
rect 64 293 68 294
rect 64 291 65 293
rect 67 291 68 293
rect 108 292 109 294
rect 111 292 112 294
rect 108 291 112 292
rect 145 293 149 294
rect 145 291 146 293
rect 148 291 149 293
rect 64 290 68 291
rect 145 290 149 291
rect 216 293 220 294
rect 216 291 217 293
rect 219 291 220 293
rect 216 290 220 291
rect 281 293 285 294
rect 281 291 282 293
rect 284 291 285 293
rect 281 290 285 291
rect 334 293 338 294
rect 402 293 406 294
rect 334 291 335 293
rect 337 291 338 293
rect 334 290 338 291
rect 369 292 373 293
rect 369 290 370 292
rect 372 290 373 292
rect 402 291 403 293
rect 405 291 406 293
rect 402 290 406 291
rect 448 293 452 294
rect 448 291 449 293
rect 451 291 452 293
rect 448 290 452 291
rect 493 293 497 294
rect 751 293 755 294
rect 493 291 494 293
rect 496 291 497 293
rect 493 290 497 291
rect 566 292 570 293
rect 566 290 567 292
rect 569 290 570 292
rect 369 289 373 290
rect 566 289 570 290
rect 631 292 635 293
rect 631 290 632 292
rect 634 290 635 292
rect 751 291 752 293
rect 754 291 755 293
rect 751 290 755 291
rect 631 289 635 290
rect 394 283 486 284
rect 394 281 395 283
rect 397 281 483 283
rect 485 281 486 283
rect 394 280 486 281
rect 227 269 333 270
rect 227 267 228 269
rect 230 267 330 269
rect 332 267 333 269
rect 227 266 333 267
rect 72 261 131 262
rect 72 259 73 261
rect 75 259 128 261
rect 130 259 131 261
rect 72 258 131 259
rect 161 261 232 262
rect 161 259 162 261
rect 164 259 229 261
rect 231 259 232 261
rect 161 258 232 259
rect 329 261 333 262
rect 329 259 330 261
rect 332 259 333 261
rect 329 258 333 259
rect 482 261 486 262
rect 482 259 483 261
rect 485 259 486 261
rect 482 258 486 259
rect 583 261 587 262
rect 583 259 584 261
rect 586 259 587 261
rect 583 258 587 259
rect 682 261 686 262
rect 682 259 683 261
rect 685 259 686 261
rect 682 258 686 259
rect 145 253 149 254
rect 500 253 504 254
rect 690 253 694 254
rect 94 252 98 253
rect 94 250 95 252
rect 97 250 98 252
rect 94 245 98 250
rect 145 251 146 253
rect 148 252 297 253
rect 148 251 294 252
rect 145 250 294 251
rect 296 250 297 252
rect 437 252 441 253
rect 437 250 438 252
rect 440 250 441 252
rect 145 249 297 250
rect 346 249 418 250
rect 346 247 347 249
rect 349 247 415 249
rect 417 247 418 249
rect 346 246 418 247
rect 437 245 441 250
rect 500 251 501 253
rect 503 252 652 253
rect 503 251 649 252
rect 500 250 649 251
rect 651 250 652 252
rect 690 251 691 253
rect 693 251 694 253
rect 690 250 694 251
rect 500 249 652 250
rect 94 244 216 245
rect 94 242 213 244
rect 215 242 216 244
rect 94 241 216 242
rect 245 244 317 245
rect 245 242 246 244
rect 248 242 314 244
rect 316 242 317 244
rect 245 241 317 242
rect 437 244 571 245
rect 437 242 568 244
rect 570 242 571 244
rect 437 241 571 242
rect 600 244 670 245
rect 600 242 601 244
rect 603 242 667 244
rect 669 242 670 244
rect 600 241 670 242
rect 236 236 587 237
rect 236 234 237 236
rect 239 234 584 236
rect 586 234 587 236
rect 236 233 587 234
rect 100 228 686 229
rect 100 226 101 228
rect 103 226 683 228
rect 685 226 686 228
rect 67 225 71 226
rect 100 225 686 226
rect 708 225 712 226
rect 67 223 68 225
rect 70 223 71 225
rect 67 222 71 223
rect 708 223 709 225
rect 711 223 712 225
rect 708 222 712 223
rect 751 225 755 226
rect 751 223 752 225
rect 754 223 755 225
rect 751 222 755 223
rect 128 220 132 221
rect 128 218 129 220
rect 131 218 132 220
rect 128 217 132 218
rect 192 220 196 221
rect 192 218 193 220
rect 195 218 196 220
rect 192 217 196 218
rect 256 220 260 221
rect 256 218 257 220
rect 259 218 260 220
rect 256 217 260 218
rect 319 220 323 221
rect 319 218 320 220
rect 322 218 323 220
rect 319 217 323 218
rect 355 220 359 221
rect 355 218 356 220
rect 358 218 359 220
rect 355 217 359 218
rect 386 220 390 221
rect 386 218 387 220
rect 389 218 390 220
rect 386 217 390 218
rect 427 220 431 221
rect 427 218 428 220
rect 430 218 431 220
rect 427 217 431 218
rect 458 220 462 221
rect 458 218 459 220
rect 461 218 462 220
rect 458 217 462 218
rect 515 220 519 221
rect 515 218 516 220
rect 518 218 519 220
rect 515 217 519 218
rect 605 220 609 221
rect 605 218 606 220
rect 608 218 609 220
rect 605 217 609 218
<< alu3 >>
rect 402 581 406 582
rect 402 579 403 581
rect 405 579 406 581
rect 107 578 111 579
rect 402 578 406 579
rect 448 581 452 582
rect 448 579 449 581
rect 451 579 452 581
rect 448 578 452 579
rect 493 581 497 582
rect 493 579 494 581
rect 496 579 497 581
rect 493 578 497 579
rect 566 581 570 582
rect 566 579 567 581
rect 569 579 570 581
rect 566 578 570 579
rect 752 578 756 579
rect 67 577 71 578
rect 67 575 68 577
rect 70 575 71 577
rect 107 576 108 578
rect 110 576 111 578
rect 107 575 111 576
rect 145 577 149 578
rect 145 575 146 577
rect 148 575 149 577
rect 67 574 71 575
rect 145 574 149 575
rect 216 577 220 578
rect 216 575 217 577
rect 219 575 220 577
rect 216 574 220 575
rect 281 577 285 578
rect 281 575 282 577
rect 284 575 285 577
rect 281 574 285 575
rect 334 577 338 578
rect 334 575 335 577
rect 337 575 338 577
rect 334 574 338 575
rect 369 577 373 578
rect 369 575 370 577
rect 372 575 373 577
rect 369 574 373 575
rect 631 577 635 578
rect 631 575 632 577
rect 634 575 635 577
rect 752 576 753 578
rect 755 576 756 578
rect 752 575 756 576
rect 631 574 635 575
rect 400 573 404 574
rect 400 571 401 573
rect 403 571 404 573
rect 167 565 171 566
rect 167 563 168 565
rect 170 563 171 565
rect 111 557 115 558
rect 111 555 112 557
rect 114 555 115 557
rect 111 549 115 555
rect 111 547 112 549
rect 114 547 115 549
rect 111 546 115 547
rect 167 549 171 563
rect 167 547 168 549
rect 170 547 171 549
rect 167 546 171 547
rect 313 565 317 566
rect 313 563 314 565
rect 316 563 317 565
rect 313 549 317 563
rect 313 547 314 549
rect 316 547 317 549
rect 313 546 317 547
rect 400 549 404 571
rect 596 573 600 574
rect 596 571 597 573
rect 599 571 600 573
rect 400 547 401 549
rect 403 547 404 549
rect 400 546 404 547
rect 483 565 487 566
rect 483 563 484 565
rect 486 563 487 565
rect 483 549 487 563
rect 483 547 484 549
rect 486 547 487 549
rect 483 546 487 547
rect 539 557 543 558
rect 539 555 540 557
rect 542 555 543 557
rect 539 549 543 555
rect 539 547 540 549
rect 542 547 543 549
rect 539 546 543 547
rect 596 549 600 571
rect 596 547 597 549
rect 599 547 600 549
rect 596 546 600 547
rect 683 565 687 566
rect 683 563 684 565
rect 686 563 687 565
rect 683 549 687 563
rect 683 547 684 549
rect 686 547 687 549
rect 683 546 687 547
rect 78 541 82 542
rect 78 539 79 541
rect 81 539 82 541
rect 78 532 82 539
rect 402 541 406 542
rect 402 539 403 541
rect 405 539 406 541
rect 78 530 79 532
rect 81 530 82 532
rect 67 509 71 510
rect 67 507 68 509
rect 70 507 71 509
rect 67 506 71 507
rect 78 486 82 530
rect 78 484 79 486
rect 81 484 82 486
rect 78 483 82 484
rect 118 532 122 533
rect 118 530 119 532
rect 121 530 122 532
rect 118 486 122 530
rect 184 532 188 533
rect 184 530 185 532
rect 187 530 188 532
rect 169 525 173 526
rect 146 524 150 525
rect 146 522 147 524
rect 149 522 150 524
rect 128 509 132 510
rect 128 507 129 509
rect 131 507 132 509
rect 128 506 132 507
rect 118 484 119 486
rect 121 484 122 486
rect 118 483 122 484
rect 99 477 103 478
rect 99 475 100 477
rect 102 475 103 477
rect 67 436 71 437
rect 67 434 68 436
rect 70 434 71 436
rect 67 433 71 434
rect 99 405 103 475
rect 107 469 111 470
rect 107 467 108 469
rect 110 467 111 469
rect 107 448 111 467
rect 146 469 150 522
rect 169 523 170 525
rect 172 523 173 525
rect 169 477 173 523
rect 184 494 188 530
rect 296 532 300 533
rect 296 530 297 532
rect 299 530 300 532
rect 236 525 240 526
rect 236 523 237 525
rect 239 523 240 525
rect 192 509 196 510
rect 192 507 193 509
rect 195 507 196 509
rect 192 506 196 507
rect 184 492 185 494
rect 187 492 188 494
rect 184 491 188 492
rect 169 475 170 477
rect 172 475 173 477
rect 169 474 173 475
rect 146 467 147 469
rect 149 467 150 469
rect 146 466 150 467
rect 208 469 212 470
rect 208 467 209 469
rect 211 467 212 469
rect 107 446 108 448
rect 110 446 111 448
rect 107 445 111 446
rect 153 461 157 462
rect 153 459 154 461
rect 156 459 157 461
rect 107 437 111 438
rect 107 435 108 437
rect 110 435 111 437
rect 107 434 111 435
rect 145 437 149 438
rect 145 435 146 437
rect 148 435 149 437
rect 145 434 149 435
rect 99 401 104 405
rect 90 396 96 397
rect 90 394 93 396
rect 95 394 96 396
rect 90 393 96 394
rect 72 381 76 382
rect 72 379 73 381
rect 75 379 76 381
rect 64 365 68 366
rect 64 363 65 365
rect 67 363 68 365
rect 64 362 68 363
rect 64 293 68 294
rect 64 291 65 293
rect 67 291 68 293
rect 64 290 68 291
rect 72 261 76 379
rect 90 349 94 393
rect 90 347 91 349
rect 93 347 94 349
rect 90 346 94 347
rect 72 259 73 261
rect 75 259 76 261
rect 72 258 76 259
rect 100 228 104 401
rect 153 396 157 459
rect 200 405 204 406
rect 200 403 201 405
rect 203 403 204 405
rect 153 394 154 396
rect 156 394 157 396
rect 153 393 157 394
rect 161 396 165 397
rect 161 394 162 396
rect 164 394 165 396
rect 152 388 156 389
rect 152 386 153 388
rect 155 386 156 388
rect 128 364 132 365
rect 128 362 129 364
rect 131 362 132 364
rect 128 361 132 362
rect 152 349 156 386
rect 152 347 153 349
rect 155 347 156 349
rect 152 346 156 347
rect 108 294 112 295
rect 108 292 109 294
rect 111 292 112 294
rect 108 291 112 292
rect 145 293 149 294
rect 145 291 146 293
rect 148 291 149 293
rect 145 290 149 291
rect 161 261 165 394
rect 200 389 204 403
rect 200 387 201 389
rect 203 387 204 389
rect 200 386 204 387
rect 184 381 188 382
rect 184 379 185 381
rect 187 379 188 381
rect 184 334 188 379
rect 192 365 196 366
rect 192 363 193 365
rect 195 363 196 365
rect 192 362 196 363
rect 184 332 185 334
rect 187 332 188 334
rect 184 331 188 332
rect 208 325 212 467
rect 227 458 231 459
rect 227 456 228 458
rect 230 456 231 458
rect 216 437 220 438
rect 216 435 217 437
rect 219 435 220 437
rect 216 434 220 435
rect 208 323 209 325
rect 211 323 212 325
rect 208 322 212 323
rect 216 293 220 294
rect 216 291 217 293
rect 219 291 220 293
rect 216 290 220 291
rect 227 269 231 456
rect 227 267 228 269
rect 230 267 231 269
rect 227 266 231 267
rect 161 259 162 261
rect 164 259 165 261
rect 161 258 165 259
rect 236 236 240 523
rect 248 525 253 526
rect 248 523 250 525
rect 252 523 253 525
rect 248 522 253 523
rect 248 477 252 522
rect 256 509 260 510
rect 256 507 257 509
rect 259 507 260 509
rect 256 506 260 507
rect 296 494 300 530
rect 362 532 366 533
rect 362 530 363 532
rect 365 530 366 532
rect 296 492 297 494
rect 299 492 300 494
rect 296 491 300 492
rect 311 525 315 526
rect 311 523 312 525
rect 314 523 315 525
rect 248 475 249 477
rect 251 475 252 477
rect 248 474 252 475
rect 297 477 301 478
rect 297 475 298 477
rect 300 475 301 477
rect 258 469 262 470
rect 258 467 259 469
rect 261 467 262 469
rect 258 461 262 467
rect 258 459 259 461
rect 261 459 262 461
rect 249 458 253 459
rect 258 458 262 459
rect 249 456 250 458
rect 252 456 253 458
rect 249 405 253 456
rect 281 437 285 438
rect 281 435 282 437
rect 284 435 285 437
rect 281 434 285 435
rect 297 413 301 475
rect 311 477 315 523
rect 334 524 338 525
rect 334 522 335 524
rect 337 522 338 524
rect 319 509 323 510
rect 319 507 320 509
rect 322 507 323 509
rect 319 506 323 507
rect 311 475 312 477
rect 314 475 315 477
rect 311 474 315 475
rect 334 469 338 522
rect 354 509 358 510
rect 354 507 355 509
rect 357 507 358 509
rect 354 506 358 507
rect 362 486 366 530
rect 402 532 406 539
rect 532 540 536 541
rect 532 538 533 540
rect 535 538 536 540
rect 402 530 403 532
rect 405 530 406 532
rect 386 509 390 510
rect 386 507 387 509
rect 389 507 390 509
rect 386 506 390 507
rect 362 484 363 486
rect 365 484 366 486
rect 362 483 366 484
rect 402 486 406 530
rect 466 532 470 533
rect 466 530 467 532
rect 469 530 470 532
rect 402 484 403 486
rect 405 484 406 486
rect 402 483 406 484
rect 419 525 423 526
rect 419 523 420 525
rect 422 523 423 525
rect 334 467 335 469
rect 337 467 338 469
rect 334 466 338 467
rect 400 469 404 470
rect 400 467 401 469
rect 403 467 404 469
rect 378 456 382 457
rect 378 454 379 456
rect 381 454 382 456
rect 334 437 338 438
rect 334 435 335 437
rect 337 435 338 437
rect 334 434 338 435
rect 369 436 373 437
rect 369 434 370 436
rect 372 434 373 436
rect 369 433 373 434
rect 297 411 298 413
rect 300 411 301 413
rect 297 410 301 411
rect 330 421 334 422
rect 330 419 331 421
rect 333 419 334 421
rect 249 403 250 405
rect 252 403 253 405
rect 249 402 253 403
rect 330 405 334 419
rect 378 421 382 454
rect 400 456 404 467
rect 400 454 401 456
rect 403 454 404 456
rect 400 453 404 454
rect 409 465 413 466
rect 409 463 410 465
rect 412 463 413 465
rect 401 436 405 437
rect 401 434 402 436
rect 404 434 405 436
rect 401 433 405 434
rect 378 419 379 421
rect 381 419 382 421
rect 378 418 382 419
rect 330 403 331 405
rect 333 403 334 405
rect 330 402 334 403
rect 358 405 362 406
rect 358 403 359 405
rect 361 403 362 405
rect 304 389 308 390
rect 304 387 305 389
rect 307 387 308 389
rect 246 381 250 382
rect 246 379 247 381
rect 249 379 250 381
rect 246 342 250 379
rect 304 380 308 387
rect 304 378 305 380
rect 307 378 308 380
rect 304 377 308 378
rect 347 388 351 389
rect 347 386 348 388
rect 350 386 351 388
rect 256 365 260 366
rect 256 363 257 365
rect 259 363 260 365
rect 256 362 260 363
rect 319 365 323 366
rect 319 363 320 365
rect 322 363 323 365
rect 319 362 323 363
rect 347 349 351 386
rect 358 380 362 403
rect 358 378 359 380
rect 361 378 362 380
rect 358 377 362 378
rect 394 381 398 382
rect 394 379 395 381
rect 397 379 398 381
rect 355 365 359 366
rect 355 363 356 365
rect 358 363 359 365
rect 355 362 359 363
rect 386 365 390 366
rect 386 363 387 365
rect 389 363 390 365
rect 386 362 390 363
rect 347 347 348 349
rect 350 347 351 349
rect 347 346 351 347
rect 246 340 247 342
rect 249 340 250 342
rect 246 339 250 340
rect 323 309 327 310
rect 323 307 324 309
rect 326 307 327 309
rect 323 301 327 307
rect 323 299 324 301
rect 326 299 327 301
rect 323 298 327 299
rect 281 293 285 294
rect 281 291 282 293
rect 284 291 285 293
rect 281 290 285 291
rect 334 293 338 294
rect 334 291 335 293
rect 337 291 338 293
rect 334 290 338 291
rect 369 292 373 293
rect 369 290 370 292
rect 372 290 373 292
rect 369 289 373 290
rect 394 283 398 379
rect 409 333 413 463
rect 419 372 423 523
rect 427 509 431 510
rect 427 507 428 509
rect 430 507 431 509
rect 427 506 431 507
rect 458 509 462 510
rect 458 507 459 509
rect 461 507 462 509
rect 458 506 462 507
rect 466 494 470 530
rect 532 532 536 538
rect 634 540 638 541
rect 634 538 635 540
rect 637 538 638 540
rect 532 530 533 532
rect 535 530 536 532
rect 466 492 467 494
rect 469 492 470 494
rect 466 491 470 492
rect 481 525 485 526
rect 481 523 482 525
rect 484 523 485 525
rect 458 485 462 486
rect 458 483 459 485
rect 461 483 462 485
rect 448 437 452 438
rect 448 435 449 437
rect 451 435 452 437
rect 448 434 452 435
rect 458 405 462 483
rect 481 477 485 523
rect 481 475 482 477
rect 484 475 485 477
rect 481 474 485 475
rect 504 524 508 525
rect 504 522 505 524
rect 507 522 508 524
rect 504 469 508 522
rect 515 509 519 510
rect 515 507 516 509
rect 518 507 519 509
rect 515 506 519 507
rect 532 486 536 530
rect 532 484 533 486
rect 535 484 536 486
rect 532 483 536 484
rect 572 532 576 533
rect 572 530 573 532
rect 575 530 576 532
rect 572 486 576 530
rect 572 484 573 486
rect 575 484 576 486
rect 572 483 576 484
rect 594 532 598 533
rect 594 530 595 532
rect 597 530 598 532
rect 594 486 598 530
rect 634 532 638 538
rect 634 530 635 532
rect 637 530 638 532
rect 605 509 609 510
rect 605 507 606 509
rect 608 507 609 509
rect 605 506 609 507
rect 594 484 595 486
rect 597 484 598 486
rect 594 483 598 484
rect 634 486 638 530
rect 700 532 704 533
rect 700 530 701 532
rect 703 530 704 532
rect 685 525 689 526
rect 634 484 635 486
rect 637 484 638 486
rect 634 483 638 484
rect 662 524 666 525
rect 662 522 663 524
rect 665 522 666 524
rect 558 477 562 478
rect 558 475 559 477
rect 561 475 562 477
rect 504 467 505 469
rect 507 467 508 469
rect 504 466 508 467
rect 539 469 543 470
rect 539 467 540 469
rect 542 467 543 469
rect 539 448 543 467
rect 539 446 540 448
rect 542 446 543 448
rect 539 445 543 446
rect 493 437 497 438
rect 493 435 494 437
rect 496 435 497 437
rect 493 434 497 435
rect 458 403 459 405
rect 461 403 462 405
rect 458 402 462 403
rect 483 413 487 414
rect 483 411 484 413
rect 486 411 487 413
rect 483 405 487 411
rect 558 413 562 475
rect 596 469 600 470
rect 596 467 597 469
rect 599 467 600 469
rect 596 456 600 467
rect 662 469 666 522
rect 685 523 686 525
rect 688 523 689 525
rect 685 477 689 523
rect 700 494 704 530
rect 708 509 712 510
rect 708 507 709 509
rect 711 507 712 509
rect 708 506 712 507
rect 752 509 756 510
rect 752 507 753 509
rect 755 507 756 509
rect 752 506 756 507
rect 700 492 701 494
rect 703 492 704 494
rect 700 491 704 492
rect 685 475 686 477
rect 688 475 689 477
rect 685 474 689 475
rect 662 467 663 469
rect 665 467 666 469
rect 662 466 666 467
rect 596 454 597 456
rect 599 454 600 456
rect 596 453 600 454
rect 653 461 657 462
rect 653 459 654 461
rect 656 459 657 461
rect 566 436 570 437
rect 566 434 567 436
rect 569 434 570 436
rect 566 433 570 434
rect 631 436 635 437
rect 631 434 632 436
rect 634 434 635 436
rect 631 433 635 434
rect 558 411 559 413
rect 561 411 562 413
rect 558 410 562 411
rect 483 403 484 405
rect 486 403 487 405
rect 483 402 487 403
rect 584 405 588 406
rect 584 403 585 405
rect 587 403 588 405
rect 419 370 420 372
rect 422 370 423 372
rect 419 369 423 370
rect 544 380 548 381
rect 544 378 545 380
rect 547 378 548 380
rect 427 364 431 365
rect 427 362 428 364
rect 430 362 431 364
rect 427 361 431 362
rect 458 364 462 365
rect 458 362 459 364
rect 461 362 462 364
rect 458 361 462 362
rect 515 364 519 365
rect 515 362 516 364
rect 518 362 519 364
rect 515 361 519 362
rect 409 331 410 333
rect 412 331 413 333
rect 409 330 413 331
rect 544 325 548 378
rect 584 372 588 403
rect 584 370 585 372
rect 587 370 588 372
rect 584 369 588 370
rect 605 365 609 366
rect 605 363 606 365
rect 608 363 609 365
rect 605 362 609 363
rect 544 323 545 325
rect 547 323 548 325
rect 653 326 657 459
rect 739 453 743 454
rect 739 451 740 453
rect 742 451 743 453
rect 683 421 687 422
rect 683 419 684 421
rect 686 419 687 421
rect 683 405 687 419
rect 683 403 684 405
rect 686 403 687 405
rect 683 402 687 403
rect 691 413 695 414
rect 691 411 692 413
rect 694 411 695 413
rect 691 397 695 411
rect 691 395 692 397
rect 694 395 695 397
rect 691 394 695 395
rect 700 381 704 382
rect 700 379 701 381
rect 703 379 704 381
rect 700 342 704 379
rect 708 365 712 366
rect 708 363 709 365
rect 711 363 712 365
rect 708 362 712 363
rect 700 340 701 342
rect 703 340 704 342
rect 700 339 704 340
rect 653 324 654 326
rect 656 324 657 326
rect 653 323 657 324
rect 739 325 743 451
rect 752 438 756 439
rect 752 436 753 438
rect 755 436 756 438
rect 752 435 756 436
rect 752 365 756 366
rect 752 363 753 365
rect 755 363 756 365
rect 752 362 756 363
rect 739 323 740 325
rect 742 323 743 325
rect 544 322 548 323
rect 739 322 743 323
rect 690 301 694 302
rect 690 299 691 301
rect 693 299 694 301
rect 402 293 406 294
rect 402 291 403 293
rect 405 291 406 293
rect 402 290 406 291
rect 448 293 452 294
rect 448 291 449 293
rect 451 291 452 293
rect 448 290 452 291
rect 493 293 497 294
rect 493 291 494 293
rect 496 291 497 293
rect 493 290 497 291
rect 566 292 570 293
rect 566 290 567 292
rect 569 290 570 292
rect 566 289 570 290
rect 631 292 635 293
rect 631 290 632 292
rect 634 290 635 292
rect 631 289 635 290
rect 394 281 395 283
rect 397 281 398 283
rect 394 280 398 281
rect 482 283 486 284
rect 482 281 483 283
rect 485 281 486 283
rect 329 269 333 270
rect 329 267 330 269
rect 332 267 333 269
rect 329 261 333 267
rect 329 259 330 261
rect 332 259 333 261
rect 329 258 333 259
rect 482 261 486 281
rect 482 259 483 261
rect 485 259 486 261
rect 482 258 486 259
rect 583 261 587 262
rect 583 259 584 261
rect 586 259 587 261
rect 236 234 237 236
rect 239 234 240 236
rect 236 233 240 234
rect 583 236 587 259
rect 583 234 584 236
rect 586 234 587 236
rect 583 233 587 234
rect 682 261 686 262
rect 682 259 683 261
rect 685 259 686 261
rect 100 226 101 228
rect 103 226 104 228
rect 67 225 71 226
rect 100 225 104 226
rect 682 228 686 259
rect 690 253 694 299
rect 751 293 755 294
rect 751 291 752 293
rect 754 291 755 293
rect 751 290 755 291
rect 690 251 691 253
rect 693 251 694 253
rect 690 250 694 251
rect 682 226 683 228
rect 685 226 686 228
rect 682 225 686 226
rect 708 225 712 226
rect 67 223 68 225
rect 70 223 71 225
rect 67 222 71 223
rect 708 223 709 225
rect 711 223 712 225
rect 708 222 712 223
rect 751 225 755 226
rect 751 223 752 225
rect 754 223 755 225
rect 751 222 755 223
rect 128 220 132 221
rect 128 218 129 220
rect 131 218 132 220
rect 128 217 132 218
rect 192 220 196 221
rect 192 218 193 220
rect 195 218 196 220
rect 192 217 196 218
rect 256 220 260 221
rect 256 218 257 220
rect 259 218 260 220
rect 256 217 260 218
rect 319 220 323 221
rect 319 218 320 220
rect 322 218 323 220
rect 319 217 323 218
rect 355 220 359 221
rect 355 218 356 220
rect 358 218 359 220
rect 355 217 359 218
rect 386 220 390 221
rect 386 218 387 220
rect 389 218 390 220
rect 386 217 390 218
rect 427 220 431 221
rect 427 218 428 220
rect 430 218 431 220
rect 427 217 431 218
rect 458 220 462 221
rect 458 218 459 220
rect 461 218 462 220
rect 458 217 462 218
rect 515 220 519 221
rect 515 218 516 220
rect 518 218 519 220
rect 515 217 519 218
rect 605 220 609 221
rect 605 218 606 220
rect 608 218 609 220
rect 605 217 609 218
<< alu4 >>
rect 48 509 52 601
rect 128 600 132 601
rect 128 598 129 600
rect 131 598 132 600
rect 48 507 49 509
rect 51 507 52 509
rect 48 365 52 507
rect 48 363 49 365
rect 51 363 52 365
rect 48 225 52 363
rect 48 223 49 225
rect 51 223 52 225
rect 48 198 52 223
rect 56 577 60 593
rect 107 592 111 593
rect 107 590 108 592
rect 110 590 111 592
rect 107 578 111 590
rect 56 575 57 577
rect 59 575 60 577
rect 56 436 60 575
rect 67 577 71 578
rect 67 575 68 577
rect 70 575 71 577
rect 67 574 71 575
rect 107 576 108 578
rect 110 576 111 578
rect 67 509 71 510
rect 67 507 68 509
rect 70 507 71 509
rect 67 506 71 507
rect 107 437 111 576
rect 56 434 57 436
rect 59 434 60 436
rect 56 293 60 434
rect 67 436 71 437
rect 67 434 68 436
rect 70 434 71 436
rect 67 433 71 434
rect 107 435 108 437
rect 110 435 111 437
rect 64 365 68 366
rect 64 363 65 365
rect 67 363 68 365
rect 64 362 68 363
rect 107 295 111 435
rect 128 509 132 598
rect 192 600 196 601
rect 192 598 193 600
rect 195 598 196 600
rect 128 507 129 509
rect 131 507 132 509
rect 128 364 132 507
rect 128 362 129 364
rect 131 362 132 364
rect 107 294 112 295
rect 56 291 57 293
rect 59 291 60 293
rect 56 207 60 291
rect 64 293 68 294
rect 64 291 65 293
rect 67 291 68 293
rect 64 290 68 291
rect 107 292 109 294
rect 111 292 112 294
rect 107 291 112 292
rect 67 225 71 226
rect 67 223 68 225
rect 70 223 71 225
rect 67 222 71 223
rect 107 210 111 291
rect 107 208 108 210
rect 110 208 111 210
rect 107 207 111 208
rect 128 220 132 362
rect 128 218 129 220
rect 131 218 132 220
rect 128 202 132 218
rect 145 592 149 593
rect 145 590 146 592
rect 148 590 149 592
rect 145 577 149 590
rect 145 575 146 577
rect 148 575 149 577
rect 145 437 149 575
rect 145 435 146 437
rect 148 435 149 437
rect 145 293 149 435
rect 145 291 146 293
rect 148 291 149 293
rect 145 210 149 291
rect 145 208 146 210
rect 148 208 149 210
rect 145 207 149 208
rect 192 509 196 598
rect 256 600 260 601
rect 256 598 257 600
rect 259 598 260 600
rect 192 507 193 509
rect 195 507 196 509
rect 192 365 196 507
rect 192 363 193 365
rect 195 363 196 365
rect 192 220 196 363
rect 192 218 193 220
rect 195 218 196 220
rect 128 200 129 202
rect 131 200 132 202
rect 128 199 132 200
rect 192 202 196 218
rect 216 592 220 593
rect 216 590 217 592
rect 219 590 220 592
rect 216 577 220 590
rect 216 575 217 577
rect 219 575 220 577
rect 216 437 220 575
rect 216 435 217 437
rect 219 435 220 437
rect 216 293 220 435
rect 216 291 217 293
rect 219 291 220 293
rect 216 210 220 291
rect 216 208 217 210
rect 219 208 220 210
rect 216 207 220 208
rect 256 509 260 598
rect 319 600 323 601
rect 319 598 320 600
rect 322 598 323 600
rect 256 507 257 509
rect 259 507 260 509
rect 256 365 260 507
rect 256 363 257 365
rect 259 363 260 365
rect 256 220 260 363
rect 256 218 257 220
rect 259 218 260 220
rect 192 200 193 202
rect 195 200 196 202
rect 192 199 196 200
rect 256 202 260 218
rect 281 592 285 593
rect 281 590 282 592
rect 284 590 285 592
rect 281 577 285 590
rect 281 575 282 577
rect 284 575 285 577
rect 281 437 285 575
rect 281 435 282 437
rect 284 435 285 437
rect 281 293 285 435
rect 281 291 282 293
rect 284 291 285 293
rect 281 210 285 291
rect 281 208 282 210
rect 284 208 285 210
rect 281 207 285 208
rect 319 509 323 598
rect 355 600 359 601
rect 355 598 356 600
rect 358 598 359 600
rect 319 507 320 509
rect 322 507 323 509
rect 319 365 323 507
rect 319 363 320 365
rect 322 363 323 365
rect 319 220 323 363
rect 319 218 320 220
rect 322 218 323 220
rect 256 200 257 202
rect 259 200 260 202
rect 256 199 260 200
rect 319 202 323 218
rect 334 592 338 593
rect 334 590 335 592
rect 337 590 338 592
rect 334 577 338 590
rect 334 575 335 577
rect 337 575 338 577
rect 334 437 338 575
rect 355 510 359 598
rect 386 600 390 601
rect 386 598 387 600
rect 389 598 390 600
rect 354 509 359 510
rect 354 507 355 509
rect 357 507 359 509
rect 354 506 359 507
rect 334 435 335 437
rect 337 435 338 437
rect 334 293 338 435
rect 334 291 335 293
rect 337 291 338 293
rect 334 210 338 291
rect 334 208 335 210
rect 337 208 338 210
rect 334 207 338 208
rect 355 365 359 506
rect 355 363 356 365
rect 358 363 359 365
rect 355 220 359 363
rect 355 218 356 220
rect 358 218 359 220
rect 319 200 320 202
rect 322 200 323 202
rect 319 199 323 200
rect 355 202 359 218
rect 369 592 373 593
rect 369 590 370 592
rect 372 590 373 592
rect 369 577 373 590
rect 369 575 370 577
rect 372 575 373 577
rect 369 436 373 575
rect 369 434 370 436
rect 372 434 373 436
rect 369 292 373 434
rect 369 290 370 292
rect 372 290 373 292
rect 369 210 373 290
rect 369 208 370 210
rect 372 208 373 210
rect 369 207 373 208
rect 386 509 390 598
rect 427 600 431 601
rect 427 598 428 600
rect 430 598 431 600
rect 386 507 387 509
rect 389 507 390 509
rect 386 365 390 507
rect 402 592 406 593
rect 402 590 403 592
rect 405 590 406 592
rect 402 581 406 590
rect 402 579 403 581
rect 405 579 406 581
rect 402 437 406 579
rect 401 436 406 437
rect 401 434 402 436
rect 404 434 406 436
rect 401 433 406 434
rect 386 363 387 365
rect 389 363 390 365
rect 386 220 390 363
rect 386 218 387 220
rect 389 218 390 220
rect 355 200 356 202
rect 358 200 359 202
rect 355 199 359 200
rect 386 202 390 218
rect 402 293 406 433
rect 402 291 403 293
rect 405 291 406 293
rect 402 210 406 291
rect 402 208 403 210
rect 405 208 406 210
rect 402 207 406 208
rect 427 509 431 598
rect 458 600 462 601
rect 458 598 459 600
rect 461 598 462 600
rect 427 507 428 509
rect 430 507 431 509
rect 427 364 431 507
rect 427 362 428 364
rect 430 362 431 364
rect 427 220 431 362
rect 427 218 428 220
rect 430 218 431 220
rect 386 200 387 202
rect 389 200 390 202
rect 386 199 390 200
rect 427 202 431 218
rect 448 592 452 593
rect 448 590 449 592
rect 451 590 452 592
rect 448 581 452 590
rect 448 579 449 581
rect 451 579 452 581
rect 448 437 452 579
rect 448 435 449 437
rect 451 435 452 437
rect 448 293 452 435
rect 448 291 449 293
rect 451 291 452 293
rect 448 210 452 291
rect 448 208 449 210
rect 451 208 452 210
rect 448 207 452 208
rect 458 509 462 598
rect 515 600 519 601
rect 515 598 516 600
rect 518 598 519 600
rect 458 507 459 509
rect 461 507 462 509
rect 458 364 462 507
rect 458 362 459 364
rect 461 362 462 364
rect 458 220 462 362
rect 458 218 459 220
rect 461 218 462 220
rect 427 200 428 202
rect 430 200 431 202
rect 427 199 431 200
rect 458 202 462 218
rect 493 592 497 593
rect 493 590 494 592
rect 496 590 497 592
rect 493 581 497 590
rect 493 579 494 581
rect 496 579 497 581
rect 493 437 497 579
rect 493 435 494 437
rect 496 435 497 437
rect 493 293 497 435
rect 493 291 494 293
rect 496 291 497 293
rect 493 210 497 291
rect 493 208 494 210
rect 496 208 497 210
rect 493 207 497 208
rect 515 509 519 598
rect 605 600 609 601
rect 605 598 606 600
rect 608 598 609 600
rect 515 507 516 509
rect 518 507 519 509
rect 515 364 519 507
rect 515 362 516 364
rect 518 362 519 364
rect 515 220 519 362
rect 515 218 516 220
rect 518 218 519 220
rect 458 200 459 202
rect 461 200 462 202
rect 458 199 462 200
rect 515 202 519 218
rect 566 592 570 593
rect 566 590 567 592
rect 569 590 570 592
rect 566 581 570 590
rect 566 579 567 581
rect 569 579 570 581
rect 566 436 570 579
rect 566 434 567 436
rect 569 434 570 436
rect 566 292 570 434
rect 566 290 567 292
rect 569 290 570 292
rect 566 210 570 290
rect 566 208 567 210
rect 569 208 570 210
rect 566 207 570 208
rect 605 509 609 598
rect 708 600 712 601
rect 708 598 709 600
rect 711 598 712 600
rect 605 507 606 509
rect 608 507 609 509
rect 605 365 609 507
rect 605 363 606 365
rect 608 363 609 365
rect 605 220 609 363
rect 605 218 606 220
rect 608 218 609 220
rect 515 200 516 202
rect 518 200 519 202
rect 515 199 519 200
rect 605 202 609 218
rect 631 592 635 593
rect 631 590 632 592
rect 634 590 635 592
rect 631 577 635 590
rect 631 575 632 577
rect 634 575 635 577
rect 631 436 635 575
rect 631 434 632 436
rect 634 434 635 436
rect 631 292 635 434
rect 631 290 632 292
rect 634 290 635 292
rect 631 210 635 290
rect 631 208 632 210
rect 634 208 635 210
rect 631 207 635 208
rect 708 509 712 598
rect 752 578 756 579
rect 752 576 753 578
rect 755 576 756 578
rect 752 575 756 576
rect 762 578 766 593
rect 762 576 763 578
rect 765 576 766 578
rect 708 507 709 509
rect 711 507 712 509
rect 708 365 712 507
rect 752 509 756 510
rect 752 507 753 509
rect 755 507 756 509
rect 752 506 756 507
rect 752 438 756 439
rect 752 436 753 438
rect 755 436 756 438
rect 752 435 756 436
rect 762 438 766 576
rect 762 436 763 438
rect 765 436 766 438
rect 708 363 709 365
rect 711 363 712 365
rect 708 225 712 363
rect 752 365 756 366
rect 752 363 753 365
rect 755 363 756 365
rect 752 362 756 363
rect 751 293 755 294
rect 751 291 752 293
rect 754 291 755 293
rect 751 290 755 291
rect 762 293 766 436
rect 762 291 763 293
rect 765 291 766 293
rect 708 223 709 225
rect 711 223 712 225
rect 605 200 606 202
rect 608 200 609 202
rect 605 199 609 200
rect 708 202 712 223
rect 751 225 755 226
rect 751 223 752 225
rect 754 223 755 225
rect 751 222 755 223
rect 762 207 766 291
rect 770 509 774 601
rect 770 507 771 509
rect 773 507 774 509
rect 770 365 774 507
rect 770 363 771 365
rect 773 363 774 365
rect 770 225 774 363
rect 770 223 771 225
rect 773 223 774 225
rect 708 200 709 202
rect 711 200 712 202
rect 708 199 712 200
rect 770 199 774 223
<< alu5 >>
rect 48 600 774 601
rect 48 598 129 600
rect 131 598 193 600
rect 195 598 257 600
rect 259 598 320 600
rect 322 598 356 600
rect 358 598 387 600
rect 389 598 428 600
rect 430 598 459 600
rect 461 598 516 600
rect 518 598 606 600
rect 608 598 709 600
rect 711 598 774 600
rect 48 597 774 598
rect 56 592 766 593
rect 56 590 108 592
rect 110 590 146 592
rect 148 590 217 592
rect 219 590 282 592
rect 284 590 335 592
rect 337 590 370 592
rect 372 590 403 592
rect 405 590 449 592
rect 451 590 494 592
rect 496 590 567 592
rect 569 590 632 592
rect 634 590 766 592
rect 56 589 766 590
rect 752 578 766 579
rect 56 577 71 578
rect 56 575 57 577
rect 59 575 68 577
rect 70 575 71 577
rect 752 576 753 578
rect 755 576 763 578
rect 765 576 766 578
rect 752 575 766 576
rect 56 574 71 575
rect 48 509 71 510
rect 48 507 49 509
rect 51 507 68 509
rect 70 507 71 509
rect 48 506 71 507
rect 752 509 774 510
rect 752 507 753 509
rect 755 507 771 509
rect 773 507 774 509
rect 752 506 774 507
rect 752 438 766 439
rect 56 436 71 437
rect 56 434 57 436
rect 59 434 68 436
rect 70 434 71 436
rect 752 436 753 438
rect 755 436 763 438
rect 765 436 766 438
rect 752 435 766 436
rect 56 433 71 434
rect 48 365 68 366
rect 48 363 49 365
rect 51 363 65 365
rect 67 363 68 365
rect 48 362 68 363
rect 752 365 774 366
rect 752 363 753 365
rect 755 363 771 365
rect 773 363 774 365
rect 752 362 774 363
rect 56 293 68 294
rect 56 291 57 293
rect 59 291 65 293
rect 67 291 68 293
rect 56 290 68 291
rect 751 293 766 294
rect 751 291 752 293
rect 754 291 763 293
rect 765 291 766 293
rect 751 290 766 291
rect 48 225 71 226
rect 48 223 49 225
rect 51 223 68 225
rect 70 223 71 225
rect 48 222 71 223
rect 751 225 774 226
rect 751 223 752 225
rect 754 223 771 225
rect 773 223 774 225
rect 751 222 774 223
rect 56 210 766 211
rect 56 208 108 210
rect 110 208 146 210
rect 148 208 217 210
rect 219 208 282 210
rect 284 208 335 210
rect 337 208 370 210
rect 372 208 403 210
rect 405 208 449 210
rect 451 208 494 210
rect 496 208 567 210
rect 569 208 632 210
rect 634 208 766 210
rect 56 207 766 208
rect 48 202 774 203
rect 48 200 129 202
rect 131 200 193 202
rect 195 200 257 202
rect 259 200 320 202
rect 322 200 356 202
rect 358 200 387 202
rect 389 200 428 202
rect 430 200 459 202
rect 461 200 516 202
rect 518 200 606 202
rect 608 200 709 202
rect 711 200 774 202
rect 48 199 774 200
<< ptie >>
rect 96 367 106 373
rect 440 371 450 373
rect 440 369 444 371
rect 446 369 450 371
rect 440 367 450 369
rect 186 359 196 361
rect 186 357 190 359
rect 192 357 196 359
rect 186 355 196 357
rect 440 359 450 361
rect 440 357 444 359
rect 446 357 450 359
rect 440 355 450 357
rect 96 227 106 229
rect 96 225 100 227
rect 102 225 106 227
rect 96 223 106 225
rect 439 227 449 229
rect 439 225 443 227
rect 445 225 449 227
rect 439 223 449 225
<< nmos >>
rect 78 521 80 534
rect 85 521 87 534
rect 98 520 100 534
rect 118 521 120 534
rect 125 521 127 534
rect 138 520 140 534
rect 159 514 161 528
rect 170 514 172 534
rect 177 514 179 534
rect 197 520 199 534
rect 207 520 209 534
rect 217 517 219 527
rect 227 514 229 527
rect 255 514 257 527
rect 265 517 267 527
rect 275 520 277 534
rect 285 520 287 534
rect 305 514 307 534
rect 312 514 314 534
rect 323 514 325 528
rect 344 520 346 534
rect 357 521 359 534
rect 364 521 366 534
rect 384 520 386 534
rect 397 521 399 534
rect 404 521 406 534
rect 425 514 427 527
rect 435 517 437 527
rect 445 520 447 534
rect 455 520 457 534
rect 475 514 477 534
rect 482 514 484 534
rect 493 514 495 528
rect 514 520 516 534
rect 527 521 529 534
rect 534 521 536 534
rect 554 520 556 534
rect 567 521 569 534
rect 574 521 576 534
rect 594 521 596 534
rect 601 521 603 534
rect 614 520 616 534
rect 634 521 636 534
rect 641 521 643 534
rect 654 520 656 534
rect 675 514 677 528
rect 686 514 688 534
rect 693 514 695 534
rect 713 520 715 534
rect 723 520 725 534
rect 733 517 735 527
rect 743 514 745 527
rect 78 482 80 495
rect 85 482 87 495
rect 98 482 100 496
rect 118 482 120 495
rect 125 482 127 495
rect 138 482 140 496
rect 159 488 161 502
rect 170 482 172 502
rect 177 482 179 502
rect 197 482 199 496
rect 207 482 209 496
rect 217 489 219 499
rect 227 489 229 502
rect 255 489 257 502
rect 265 489 267 499
rect 275 482 277 496
rect 285 482 287 496
rect 305 482 307 502
rect 312 482 314 502
rect 323 488 325 502
rect 344 482 346 496
rect 357 482 359 495
rect 364 482 366 495
rect 384 482 386 496
rect 397 482 399 495
rect 404 482 406 495
rect 425 489 427 502
rect 435 489 437 499
rect 445 482 447 496
rect 455 482 457 496
rect 475 482 477 502
rect 482 482 484 502
rect 493 488 495 502
rect 514 482 516 496
rect 527 482 529 495
rect 534 482 536 495
rect 554 482 556 496
rect 567 482 569 495
rect 574 482 576 495
rect 594 482 596 495
rect 601 482 603 495
rect 614 482 616 496
rect 634 482 636 495
rect 641 482 643 495
rect 654 482 656 496
rect 675 488 677 502
rect 686 482 688 502
rect 693 482 695 502
rect 713 482 715 496
rect 723 482 725 496
rect 733 489 735 499
rect 743 489 745 502
rect 78 376 80 390
rect 88 377 90 385
rect 98 379 100 387
rect 119 370 121 384
rect 130 370 132 390
rect 137 370 139 390
rect 157 376 159 390
rect 167 376 169 390
rect 177 373 179 383
rect 187 370 189 383
rect 220 370 222 384
rect 231 370 233 390
rect 238 370 240 390
rect 258 376 260 390
rect 268 376 270 390
rect 278 373 280 383
rect 288 370 290 383
rect 322 370 324 384
rect 333 370 335 390
rect 340 370 342 390
rect 360 376 362 390
rect 370 376 372 390
rect 380 373 382 383
rect 390 370 392 383
rect 422 376 424 390
rect 432 377 434 385
rect 442 379 444 387
rect 475 370 477 384
rect 486 370 488 390
rect 493 370 495 390
rect 513 376 515 390
rect 523 376 525 390
rect 533 373 535 383
rect 543 370 545 383
rect 576 370 578 384
rect 587 370 589 390
rect 594 370 596 390
rect 614 376 616 390
rect 624 376 626 390
rect 634 373 636 383
rect 644 370 646 383
rect 675 370 677 384
rect 686 370 688 390
rect 693 370 695 390
rect 713 376 715 390
rect 723 376 725 390
rect 733 373 735 383
rect 743 370 745 383
rect 80 344 82 358
rect 91 338 93 358
rect 98 338 100 358
rect 118 338 120 352
rect 128 338 130 352
rect 138 345 140 355
rect 148 345 150 358
rect 168 338 170 352
rect 178 343 180 351
rect 188 341 190 349
rect 221 344 223 358
rect 232 338 234 358
rect 239 338 241 358
rect 259 338 261 352
rect 269 338 271 352
rect 279 345 281 355
rect 289 345 291 358
rect 321 345 323 358
rect 331 345 333 355
rect 341 338 343 352
rect 351 338 353 352
rect 371 338 373 358
rect 378 338 380 358
rect 389 344 391 358
rect 422 338 424 352
rect 432 343 434 351
rect 442 341 444 349
rect 475 344 477 358
rect 486 338 488 358
rect 493 338 495 358
rect 513 338 515 352
rect 523 338 525 352
rect 533 345 535 355
rect 543 345 545 358
rect 576 344 578 358
rect 587 338 589 358
rect 594 338 596 358
rect 614 338 616 352
rect 624 338 626 352
rect 634 345 636 355
rect 644 345 646 358
rect 675 344 677 358
rect 686 338 688 358
rect 693 338 695 358
rect 713 338 715 352
rect 723 338 725 352
rect 733 345 735 355
rect 743 345 745 358
rect 78 232 80 246
rect 88 233 90 241
rect 98 235 100 243
rect 119 226 121 240
rect 130 226 132 246
rect 137 226 139 246
rect 157 232 159 246
rect 167 232 169 246
rect 177 229 179 239
rect 187 226 189 239
rect 220 226 222 240
rect 231 226 233 246
rect 238 226 240 246
rect 258 232 260 246
rect 268 232 270 246
rect 278 229 280 239
rect 288 226 290 239
rect 321 226 323 240
rect 332 226 334 246
rect 339 226 341 246
rect 359 232 361 246
rect 369 232 371 246
rect 379 229 381 239
rect 389 226 391 239
rect 421 232 423 246
rect 431 233 433 241
rect 441 235 443 243
rect 474 226 476 240
rect 485 226 487 246
rect 492 226 494 246
rect 512 232 514 246
rect 522 232 524 246
rect 532 229 534 239
rect 542 226 544 239
rect 575 226 577 240
rect 586 226 588 246
rect 593 226 595 246
rect 613 232 615 246
rect 623 232 625 246
rect 633 229 635 239
rect 643 226 645 239
rect 674 226 676 240
rect 685 226 687 246
rect 692 226 694 246
rect 712 232 714 246
rect 722 232 724 246
rect 732 229 734 239
rect 742 226 744 239
<< pmos >>
rect 78 555 80 574
rect 88 555 90 574
rect 98 546 100 574
rect 118 555 120 574
rect 128 555 130 574
rect 138 546 140 574
rect 159 546 161 574
rect 169 546 171 574
rect 179 546 181 574
rect 197 546 199 571
rect 204 546 206 571
rect 214 549 216 562
rect 227 549 229 574
rect 255 549 257 574
rect 268 549 270 562
rect 278 546 280 571
rect 285 546 287 571
rect 303 546 305 574
rect 313 546 315 574
rect 323 546 325 574
rect 344 546 346 574
rect 354 555 356 574
rect 364 555 366 574
rect 384 546 386 574
rect 394 555 396 574
rect 404 555 406 574
rect 425 549 427 574
rect 438 549 440 562
rect 448 546 450 571
rect 455 546 457 571
rect 473 546 475 574
rect 483 546 485 574
rect 493 546 495 574
rect 514 546 516 574
rect 524 555 526 574
rect 534 555 536 574
rect 554 546 556 574
rect 564 555 566 574
rect 574 555 576 574
rect 594 555 596 574
rect 604 555 606 574
rect 614 546 616 574
rect 634 555 636 574
rect 644 555 646 574
rect 654 546 656 574
rect 675 546 677 574
rect 685 546 687 574
rect 695 546 697 574
rect 713 546 715 571
rect 720 546 722 571
rect 730 549 732 562
rect 743 549 745 574
rect 78 442 80 461
rect 88 442 90 461
rect 98 442 100 470
rect 118 442 120 461
rect 128 442 130 461
rect 138 442 140 470
rect 159 442 161 470
rect 169 442 171 470
rect 179 442 181 470
rect 197 445 199 470
rect 204 445 206 470
rect 214 454 216 467
rect 227 442 229 467
rect 255 442 257 467
rect 268 454 270 467
rect 278 445 280 470
rect 285 445 287 470
rect 303 442 305 470
rect 313 442 315 470
rect 323 442 325 470
rect 344 442 346 470
rect 354 442 356 461
rect 364 442 366 461
rect 384 442 386 470
rect 394 442 396 461
rect 404 442 406 461
rect 425 442 427 467
rect 438 454 440 467
rect 448 445 450 470
rect 455 445 457 470
rect 473 442 475 470
rect 483 442 485 470
rect 493 442 495 470
rect 514 442 516 470
rect 524 442 526 461
rect 534 442 536 461
rect 554 442 556 470
rect 564 442 566 461
rect 574 442 576 461
rect 594 442 596 461
rect 604 442 606 461
rect 614 442 616 470
rect 634 442 636 461
rect 644 442 646 461
rect 654 442 656 470
rect 675 442 677 470
rect 685 442 687 470
rect 695 442 697 470
rect 713 445 715 470
rect 720 445 722 470
rect 730 454 732 467
rect 743 442 745 467
rect 78 402 80 430
rect 91 402 93 430
rect 98 402 100 430
rect 119 402 121 430
rect 129 402 131 430
rect 139 402 141 430
rect 157 402 159 427
rect 164 402 166 427
rect 174 405 176 418
rect 187 405 189 430
rect 220 402 222 430
rect 230 402 232 430
rect 240 402 242 430
rect 258 402 260 427
rect 265 402 267 427
rect 275 405 277 418
rect 288 405 290 430
rect 322 402 324 430
rect 332 402 334 430
rect 342 402 344 430
rect 360 402 362 427
rect 367 402 369 427
rect 377 405 379 418
rect 390 405 392 430
rect 422 402 424 430
rect 435 402 437 430
rect 442 402 444 430
rect 475 402 477 430
rect 485 402 487 430
rect 495 402 497 430
rect 513 402 515 427
rect 520 402 522 427
rect 530 405 532 418
rect 543 405 545 430
rect 576 402 578 430
rect 586 402 588 430
rect 596 402 598 430
rect 614 402 616 427
rect 621 402 623 427
rect 631 405 633 418
rect 644 405 646 430
rect 675 402 677 430
rect 685 402 687 430
rect 695 402 697 430
rect 713 402 715 427
rect 720 402 722 427
rect 730 405 732 418
rect 743 405 745 430
rect 80 298 82 326
rect 90 298 92 326
rect 100 298 102 326
rect 118 301 120 326
rect 125 301 127 326
rect 135 310 137 323
rect 148 298 150 323
rect 168 298 170 326
rect 181 298 183 326
rect 188 298 190 326
rect 221 298 223 326
rect 231 298 233 326
rect 241 298 243 326
rect 259 301 261 326
rect 266 301 268 326
rect 276 310 278 323
rect 289 298 291 323
rect 321 298 323 323
rect 334 310 336 323
rect 344 301 346 326
rect 351 301 353 326
rect 369 298 371 326
rect 379 298 381 326
rect 389 298 391 326
rect 422 298 424 326
rect 435 298 437 326
rect 442 298 444 326
rect 475 298 477 326
rect 485 298 487 326
rect 495 298 497 326
rect 513 301 515 326
rect 520 301 522 326
rect 530 310 532 323
rect 543 298 545 323
rect 576 298 578 326
rect 586 298 588 326
rect 596 298 598 326
rect 614 301 616 326
rect 621 301 623 326
rect 631 310 633 323
rect 644 298 646 323
rect 675 298 677 326
rect 685 298 687 326
rect 695 298 697 326
rect 713 301 715 326
rect 720 301 722 326
rect 730 310 732 323
rect 743 298 745 323
rect 78 258 80 286
rect 91 258 93 286
rect 98 258 100 286
rect 119 258 121 286
rect 129 258 131 286
rect 139 258 141 286
rect 157 258 159 283
rect 164 258 166 283
rect 174 261 176 274
rect 187 261 189 286
rect 220 258 222 286
rect 230 258 232 286
rect 240 258 242 286
rect 258 258 260 283
rect 265 258 267 283
rect 275 261 277 274
rect 288 261 290 286
rect 321 258 323 286
rect 331 258 333 286
rect 341 258 343 286
rect 359 258 361 283
rect 366 258 368 283
rect 376 261 378 274
rect 389 261 391 286
rect 421 258 423 286
rect 434 258 436 286
rect 441 258 443 286
rect 474 258 476 286
rect 484 258 486 286
rect 494 258 496 286
rect 512 258 514 283
rect 519 258 521 283
rect 529 261 531 274
rect 542 261 544 286
rect 575 258 577 286
rect 585 258 587 286
rect 595 258 597 286
rect 613 258 615 283
rect 620 258 622 283
rect 630 261 632 274
rect 643 261 645 286
rect 674 258 676 286
rect 684 258 686 286
rect 694 258 696 286
rect 712 258 714 283
rect 719 258 721 283
rect 729 261 731 274
rect 742 261 744 286
<< polyct0 >>
rect 96 539 98 541
rect 136 539 138 541
rect 159 539 161 541
rect 169 539 171 541
rect 219 542 221 544
rect 225 532 227 534
rect 263 542 265 544
rect 257 532 259 534
rect 313 539 315 541
rect 323 539 325 541
rect 346 539 348 541
rect 386 539 388 541
rect 433 542 435 544
rect 427 532 429 534
rect 483 539 485 541
rect 493 539 495 541
rect 516 539 518 541
rect 556 539 558 541
rect 612 539 614 541
rect 652 539 654 541
rect 675 539 677 541
rect 685 539 687 541
rect 735 542 737 544
rect 741 532 743 534
rect 96 475 98 477
rect 136 475 138 477
rect 159 475 161 477
rect 169 475 171 477
rect 225 482 227 484
rect 219 472 221 474
rect 257 482 259 484
rect 263 472 265 474
rect 427 482 429 484
rect 313 475 315 477
rect 323 475 325 477
rect 346 475 348 477
rect 386 475 388 477
rect 433 472 435 474
rect 483 475 485 477
rect 493 475 495 477
rect 516 475 518 477
rect 556 475 558 477
rect 612 475 614 477
rect 652 475 654 477
rect 675 475 677 477
rect 685 475 687 477
rect 741 482 743 484
rect 735 472 737 474
rect 80 395 82 397
rect 119 395 121 397
rect 129 395 131 397
rect 179 398 181 400
rect 220 395 222 397
rect 230 395 232 397
rect 185 388 187 390
rect 280 398 282 400
rect 322 395 324 397
rect 332 395 334 397
rect 286 388 288 390
rect 382 398 384 400
rect 424 395 426 397
rect 475 395 477 397
rect 485 395 487 397
rect 388 388 390 390
rect 535 398 537 400
rect 576 395 578 397
rect 586 395 588 397
rect 541 388 543 390
rect 636 398 638 400
rect 675 395 677 397
rect 685 395 687 397
rect 642 388 644 390
rect 735 398 737 400
rect 741 388 743 390
rect 80 331 82 333
rect 90 331 92 333
rect 146 338 148 340
rect 140 328 142 330
rect 170 331 172 333
rect 221 331 223 333
rect 231 331 233 333
rect 287 338 289 340
rect 281 328 283 330
rect 323 338 325 340
rect 329 328 331 330
rect 379 331 381 333
rect 389 331 391 333
rect 424 331 426 333
rect 475 331 477 333
rect 485 331 487 333
rect 541 338 543 340
rect 535 328 537 330
rect 576 331 578 333
rect 586 331 588 333
rect 642 338 644 340
rect 636 328 638 330
rect 675 331 677 333
rect 685 331 687 333
rect 741 338 743 340
rect 735 328 737 330
rect 80 251 82 253
rect 119 251 121 253
rect 129 251 131 253
rect 179 254 181 256
rect 220 251 222 253
rect 230 251 232 253
rect 185 244 187 246
rect 280 254 282 256
rect 321 251 323 253
rect 331 251 333 253
rect 286 244 288 246
rect 381 254 383 256
rect 423 251 425 253
rect 474 251 476 253
rect 484 251 486 253
rect 387 244 389 246
rect 534 254 536 256
rect 575 251 577 253
rect 585 251 587 253
rect 540 244 542 246
rect 635 254 637 256
rect 674 251 676 253
rect 684 251 686 253
rect 641 244 643 246
rect 734 254 736 256
rect 740 244 742 246
<< polyct1 >>
rect 76 547 78 549
rect 116 547 118 549
rect 86 539 88 541
rect 126 539 128 541
rect 179 539 181 541
rect 186 539 188 541
rect 205 539 207 541
rect 366 547 368 549
rect 277 539 279 541
rect 296 539 298 541
rect 303 539 305 541
rect 356 539 358 541
rect 406 547 408 549
rect 396 539 398 541
rect 536 547 538 549
rect 447 539 449 541
rect 466 539 468 541
rect 473 539 475 541
rect 526 539 528 541
rect 576 547 578 549
rect 592 547 594 549
rect 566 539 568 541
rect 632 547 634 549
rect 602 539 604 541
rect 642 539 644 541
rect 695 539 697 541
rect 702 539 704 541
rect 721 539 723 541
rect 86 475 88 477
rect 76 467 78 469
rect 126 475 128 477
rect 179 475 181 477
rect 186 475 188 477
rect 205 475 207 477
rect 116 467 118 469
rect 277 475 279 477
rect 296 475 298 477
rect 303 475 305 477
rect 356 475 358 477
rect 396 475 398 477
rect 366 467 368 469
rect 406 467 408 469
rect 447 475 449 477
rect 466 475 468 477
rect 473 475 475 477
rect 526 475 528 477
rect 566 475 568 477
rect 536 467 538 469
rect 602 475 604 477
rect 576 467 578 469
rect 592 467 594 469
rect 642 475 644 477
rect 695 475 697 477
rect 702 475 704 477
rect 721 475 723 477
rect 632 467 634 469
rect 90 395 92 397
rect 103 395 105 397
rect 139 395 141 397
rect 146 395 148 397
rect 165 395 167 397
rect 240 395 242 397
rect 247 395 249 397
rect 266 395 268 397
rect 342 395 344 397
rect 349 395 351 397
rect 368 395 370 397
rect 434 395 436 397
rect 447 395 449 397
rect 495 395 497 397
rect 502 395 504 397
rect 521 395 523 397
rect 596 395 598 397
rect 603 395 605 397
rect 622 395 624 397
rect 695 395 697 397
rect 702 395 704 397
rect 721 395 723 397
rect 100 331 102 333
rect 107 331 109 333
rect 126 331 128 333
rect 180 331 182 333
rect 193 331 195 333
rect 241 331 243 333
rect 248 331 250 333
rect 267 331 269 333
rect 343 331 345 333
rect 362 331 364 333
rect 369 331 371 333
rect 434 331 436 333
rect 447 331 449 333
rect 495 331 497 333
rect 502 331 504 333
rect 521 331 523 333
rect 596 331 598 333
rect 603 331 605 333
rect 622 331 624 333
rect 695 331 697 333
rect 702 331 704 333
rect 721 331 723 333
rect 90 251 92 253
rect 103 251 105 253
rect 139 251 141 253
rect 146 251 148 253
rect 165 251 167 253
rect 240 251 242 253
rect 247 251 249 253
rect 266 251 268 253
rect 341 251 343 253
rect 348 251 350 253
rect 367 251 369 253
rect 433 251 435 253
rect 446 251 448 253
rect 494 251 496 253
rect 501 251 503 253
rect 520 251 522 253
rect 595 251 597 253
rect 602 251 604 253
rect 621 251 623 253
rect 694 251 696 253
rect 701 251 703 253
rect 720 251 722 253
<< ndifct0 >>
rect 73 523 75 525
rect 113 523 115 525
rect 165 516 167 518
rect 192 530 194 532
rect 182 523 184 525
rect 192 523 194 525
rect 202 530 204 532
rect 212 522 214 524
rect 222 519 224 521
rect 260 519 262 521
rect 270 522 272 524
rect 280 530 282 532
rect 290 530 292 532
rect 290 523 292 525
rect 300 523 302 525
rect 317 516 319 518
rect 369 523 371 525
rect 409 523 411 525
rect 430 519 432 521
rect 440 522 442 524
rect 450 530 452 532
rect 460 530 462 532
rect 460 523 462 525
rect 470 523 472 525
rect 487 516 489 518
rect 539 523 541 525
rect 579 523 581 525
rect 589 523 591 525
rect 629 523 631 525
rect 681 516 683 518
rect 708 530 710 532
rect 698 523 700 525
rect 708 523 710 525
rect 718 530 720 532
rect 728 522 730 524
rect 738 519 740 521
rect 73 491 75 493
rect 113 491 115 493
rect 165 498 167 500
rect 182 491 184 493
rect 192 491 194 493
rect 192 484 194 486
rect 202 484 204 486
rect 212 492 214 494
rect 222 495 224 497
rect 260 495 262 497
rect 270 492 272 494
rect 280 484 282 486
rect 290 491 292 493
rect 300 491 302 493
rect 290 484 292 486
rect 317 498 319 500
rect 369 491 371 493
rect 409 491 411 493
rect 430 495 432 497
rect 440 492 442 494
rect 450 484 452 486
rect 460 491 462 493
rect 470 491 472 493
rect 460 484 462 486
rect 487 498 489 500
rect 539 491 541 493
rect 579 491 581 493
rect 589 491 591 493
rect 629 491 631 493
rect 681 498 683 500
rect 698 491 700 493
rect 708 491 710 493
rect 708 484 710 486
rect 718 484 720 486
rect 728 492 730 494
rect 738 495 740 497
rect 83 379 85 381
rect 93 381 95 383
rect 103 381 105 383
rect 125 372 127 374
rect 152 386 154 388
rect 142 379 144 381
rect 152 379 154 381
rect 162 386 164 388
rect 172 378 174 380
rect 182 375 184 377
rect 226 372 228 374
rect 253 386 255 388
rect 243 379 245 381
rect 253 379 255 381
rect 263 386 265 388
rect 273 378 275 380
rect 283 375 285 377
rect 328 372 330 374
rect 355 386 357 388
rect 345 379 347 381
rect 355 379 357 381
rect 365 386 367 388
rect 375 378 377 380
rect 385 375 387 377
rect 427 379 429 381
rect 437 381 439 383
rect 447 381 449 383
rect 481 372 483 374
rect 508 386 510 388
rect 498 379 500 381
rect 508 379 510 381
rect 518 386 520 388
rect 528 378 530 380
rect 538 375 540 377
rect 582 372 584 374
rect 609 386 611 388
rect 599 379 601 381
rect 609 379 611 381
rect 619 386 621 388
rect 629 378 631 380
rect 639 375 641 377
rect 681 372 683 374
rect 708 386 710 388
rect 698 379 700 381
rect 708 379 710 381
rect 718 386 720 388
rect 728 378 730 380
rect 738 375 740 377
rect 86 354 88 356
rect 103 347 105 349
rect 113 347 115 349
rect 113 340 115 342
rect 123 340 125 342
rect 133 348 135 350
rect 143 351 145 353
rect 173 347 175 349
rect 183 345 185 347
rect 193 345 195 347
rect 227 354 229 356
rect 244 347 246 349
rect 254 347 256 349
rect 254 340 256 342
rect 264 340 266 342
rect 274 348 276 350
rect 284 351 286 353
rect 326 351 328 353
rect 336 348 338 350
rect 346 340 348 342
rect 356 347 358 349
rect 366 347 368 349
rect 356 340 358 342
rect 383 354 385 356
rect 427 347 429 349
rect 437 345 439 347
rect 447 345 449 347
rect 481 354 483 356
rect 498 347 500 349
rect 508 347 510 349
rect 508 340 510 342
rect 518 340 520 342
rect 528 348 530 350
rect 538 351 540 353
rect 582 354 584 356
rect 599 347 601 349
rect 609 347 611 349
rect 609 340 611 342
rect 619 340 621 342
rect 629 348 631 350
rect 639 351 641 353
rect 681 354 683 356
rect 698 347 700 349
rect 708 347 710 349
rect 708 340 710 342
rect 718 340 720 342
rect 728 348 730 350
rect 738 351 740 353
rect 83 235 85 237
rect 93 237 95 239
rect 103 237 105 239
rect 125 228 127 230
rect 152 242 154 244
rect 142 235 144 237
rect 152 235 154 237
rect 162 242 164 244
rect 172 234 174 236
rect 182 231 184 233
rect 226 228 228 230
rect 253 242 255 244
rect 243 235 245 237
rect 253 235 255 237
rect 263 242 265 244
rect 273 234 275 236
rect 283 231 285 233
rect 327 228 329 230
rect 354 242 356 244
rect 344 235 346 237
rect 354 235 356 237
rect 364 242 366 244
rect 374 234 376 236
rect 384 231 386 233
rect 426 235 428 237
rect 436 237 438 239
rect 446 237 448 239
rect 480 228 482 230
rect 507 242 509 244
rect 497 235 499 237
rect 507 235 509 237
rect 517 242 519 244
rect 527 234 529 236
rect 537 231 539 233
rect 581 228 583 230
rect 608 242 610 244
rect 598 235 600 237
rect 608 235 610 237
rect 618 242 620 244
rect 628 234 630 236
rect 638 231 640 233
rect 680 228 682 230
rect 707 242 709 244
rect 697 235 699 237
rect 707 235 709 237
rect 717 242 719 244
rect 727 234 729 236
rect 737 231 739 233
<< ndifct1 >>
rect 103 530 105 532
rect 103 522 105 524
rect 143 530 145 532
rect 143 522 145 524
rect 154 523 156 525
rect 92 513 94 515
rect 132 513 134 515
rect 232 523 234 525
rect 250 523 252 525
rect 339 530 341 532
rect 328 523 330 525
rect 339 522 341 524
rect 379 530 381 532
rect 379 522 381 524
rect 420 523 422 525
rect 350 513 352 515
rect 390 513 392 515
rect 509 530 511 532
rect 498 523 500 525
rect 509 522 511 524
rect 549 530 551 532
rect 549 522 551 524
rect 619 530 621 532
rect 619 522 621 524
rect 520 513 522 515
rect 560 513 562 515
rect 659 530 661 532
rect 659 522 661 524
rect 670 523 672 525
rect 608 513 610 515
rect 648 513 650 515
rect 748 523 750 525
rect 92 501 94 503
rect 132 501 134 503
rect 103 492 105 494
rect 103 484 105 486
rect 143 492 145 494
rect 154 491 156 493
rect 143 484 145 486
rect 232 491 234 493
rect 250 491 252 493
rect 350 501 352 503
rect 390 501 392 503
rect 328 491 330 493
rect 339 492 341 494
rect 339 484 341 486
rect 379 492 381 494
rect 379 484 381 486
rect 420 491 422 493
rect 520 501 522 503
rect 560 501 562 503
rect 498 491 500 493
rect 509 492 511 494
rect 509 484 511 486
rect 608 501 610 503
rect 648 501 650 503
rect 549 492 551 494
rect 549 484 551 486
rect 619 492 621 494
rect 619 484 621 486
rect 659 492 661 494
rect 670 491 672 493
rect 659 484 661 486
rect 748 491 750 493
rect 73 386 75 388
rect 73 379 75 381
rect 114 379 116 381
rect 192 379 194 381
rect 215 379 217 381
rect 293 379 295 381
rect 317 379 319 381
rect 417 386 419 388
rect 395 379 397 381
rect 417 379 419 381
rect 470 379 472 381
rect 548 379 550 381
rect 571 379 573 381
rect 649 379 651 381
rect 670 379 672 381
rect 748 379 750 381
rect 75 347 77 349
rect 153 347 155 349
rect 163 347 165 349
rect 163 340 165 342
rect 216 347 218 349
rect 294 347 296 349
rect 316 347 318 349
rect 394 347 396 349
rect 417 347 419 349
rect 417 340 419 342
rect 470 347 472 349
rect 548 347 550 349
rect 571 347 573 349
rect 649 347 651 349
rect 670 347 672 349
rect 748 347 750 349
rect 73 242 75 244
rect 73 235 75 237
rect 114 235 116 237
rect 192 235 194 237
rect 215 235 217 237
rect 293 235 295 237
rect 316 235 318 237
rect 416 242 418 244
rect 394 235 396 237
rect 416 235 418 237
rect 469 235 471 237
rect 547 235 549 237
rect 570 235 572 237
rect 648 235 650 237
rect 669 235 671 237
rect 747 235 749 237
<< ptiect1 >>
rect 444 369 446 371
rect 190 357 192 359
rect 444 357 446 359
rect 100 225 102 227
rect 443 225 445 227
<< pdifct0 >>
rect 73 570 75 572
rect 73 563 75 565
rect 83 564 85 566
rect 83 557 85 559
rect 93 570 95 572
rect 93 563 95 565
rect 113 570 115 572
rect 113 563 115 565
rect 123 564 125 566
rect 123 557 125 559
rect 133 570 135 572
rect 133 563 135 565
rect 164 570 166 572
rect 164 563 166 565
rect 174 562 176 564
rect 174 555 176 557
rect 186 570 188 572
rect 186 563 188 565
rect 221 570 223 572
rect 209 551 211 553
rect 261 570 263 572
rect 273 551 275 553
rect 296 570 298 572
rect 296 563 298 565
rect 308 562 310 564
rect 308 555 310 557
rect 318 570 320 572
rect 318 563 320 565
rect 349 570 351 572
rect 349 563 351 565
rect 359 564 361 566
rect 359 557 361 559
rect 369 570 371 572
rect 369 563 371 565
rect 389 570 391 572
rect 389 563 391 565
rect 399 564 401 566
rect 399 557 401 559
rect 409 570 411 572
rect 409 563 411 565
rect 431 570 433 572
rect 443 551 445 553
rect 466 570 468 572
rect 466 563 468 565
rect 478 562 480 564
rect 478 555 480 557
rect 488 570 490 572
rect 488 563 490 565
rect 519 570 521 572
rect 519 563 521 565
rect 529 564 531 566
rect 529 557 531 559
rect 539 570 541 572
rect 539 563 541 565
rect 559 570 561 572
rect 559 563 561 565
rect 569 564 571 566
rect 569 557 571 559
rect 579 570 581 572
rect 579 563 581 565
rect 589 570 591 572
rect 589 563 591 565
rect 599 564 601 566
rect 599 557 601 559
rect 609 570 611 572
rect 609 563 611 565
rect 629 570 631 572
rect 629 563 631 565
rect 639 564 641 566
rect 639 557 641 559
rect 649 570 651 572
rect 649 563 651 565
rect 680 570 682 572
rect 680 563 682 565
rect 690 562 692 564
rect 690 555 692 557
rect 702 570 704 572
rect 702 563 704 565
rect 737 570 739 572
rect 725 551 727 553
rect 73 451 75 453
rect 73 444 75 446
rect 83 457 85 459
rect 83 450 85 452
rect 93 451 95 453
rect 93 444 95 446
rect 113 451 115 453
rect 113 444 115 446
rect 123 457 125 459
rect 123 450 125 452
rect 133 451 135 453
rect 133 444 135 446
rect 164 451 166 453
rect 164 444 166 446
rect 174 459 176 461
rect 174 452 176 454
rect 186 451 188 453
rect 186 444 188 446
rect 209 463 211 465
rect 221 444 223 446
rect 273 463 275 465
rect 261 444 263 446
rect 296 451 298 453
rect 296 444 298 446
rect 308 459 310 461
rect 308 452 310 454
rect 318 451 320 453
rect 318 444 320 446
rect 349 451 351 453
rect 349 444 351 446
rect 359 457 361 459
rect 359 450 361 452
rect 369 451 371 453
rect 369 444 371 446
rect 389 451 391 453
rect 389 444 391 446
rect 399 457 401 459
rect 399 450 401 452
rect 409 451 411 453
rect 409 444 411 446
rect 443 463 445 465
rect 431 444 433 446
rect 466 451 468 453
rect 466 444 468 446
rect 478 459 480 461
rect 478 452 480 454
rect 488 451 490 453
rect 488 444 490 446
rect 519 451 521 453
rect 519 444 521 446
rect 529 457 531 459
rect 529 450 531 452
rect 539 451 541 453
rect 539 444 541 446
rect 559 451 561 453
rect 559 444 561 446
rect 569 457 571 459
rect 569 450 571 452
rect 579 451 581 453
rect 579 444 581 446
rect 589 451 591 453
rect 589 444 591 446
rect 599 457 601 459
rect 599 450 601 452
rect 609 451 611 453
rect 609 444 611 446
rect 629 451 631 453
rect 629 444 631 446
rect 639 457 641 459
rect 639 450 641 452
rect 649 451 651 453
rect 649 444 651 446
rect 680 451 682 453
rect 680 444 682 446
rect 690 459 692 461
rect 690 452 692 454
rect 702 451 704 453
rect 702 444 704 446
rect 725 463 727 465
rect 737 444 739 446
rect 103 420 105 422
rect 124 426 126 428
rect 124 419 126 421
rect 134 418 136 420
rect 134 411 136 413
rect 146 426 148 428
rect 146 419 148 421
rect 181 426 183 428
rect 169 407 171 409
rect 225 426 227 428
rect 225 419 227 421
rect 235 418 237 420
rect 235 411 237 413
rect 247 426 249 428
rect 247 419 249 421
rect 282 426 284 428
rect 270 407 272 409
rect 327 426 329 428
rect 327 419 329 421
rect 337 418 339 420
rect 337 411 339 413
rect 349 426 351 428
rect 349 419 351 421
rect 384 426 386 428
rect 372 407 374 409
rect 447 420 449 422
rect 480 426 482 428
rect 480 419 482 421
rect 490 418 492 420
rect 490 411 492 413
rect 502 426 504 428
rect 502 419 504 421
rect 537 426 539 428
rect 525 407 527 409
rect 581 426 583 428
rect 581 419 583 421
rect 591 418 593 420
rect 591 411 593 413
rect 603 426 605 428
rect 603 419 605 421
rect 638 426 640 428
rect 626 407 628 409
rect 680 426 682 428
rect 680 419 682 421
rect 690 418 692 420
rect 690 411 692 413
rect 702 426 704 428
rect 702 419 704 421
rect 737 426 739 428
rect 725 407 727 409
rect 85 307 87 309
rect 85 300 87 302
rect 95 315 97 317
rect 95 308 97 310
rect 107 307 109 309
rect 107 300 109 302
rect 130 319 132 321
rect 142 300 144 302
rect 193 306 195 308
rect 226 307 228 309
rect 226 300 228 302
rect 236 315 238 317
rect 236 308 238 310
rect 248 307 250 309
rect 248 300 250 302
rect 271 319 273 321
rect 283 300 285 302
rect 339 319 341 321
rect 327 300 329 302
rect 362 307 364 309
rect 362 300 364 302
rect 374 315 376 317
rect 374 308 376 310
rect 384 307 386 309
rect 384 300 386 302
rect 447 306 449 308
rect 480 307 482 309
rect 480 300 482 302
rect 490 315 492 317
rect 490 308 492 310
rect 502 307 504 309
rect 502 300 504 302
rect 525 319 527 321
rect 537 300 539 302
rect 581 307 583 309
rect 581 300 583 302
rect 591 315 593 317
rect 591 308 593 310
rect 603 307 605 309
rect 603 300 605 302
rect 626 319 628 321
rect 638 300 640 302
rect 680 307 682 309
rect 680 300 682 302
rect 690 315 692 317
rect 690 308 692 310
rect 702 307 704 309
rect 702 300 704 302
rect 725 319 727 321
rect 737 300 739 302
rect 103 276 105 278
rect 124 282 126 284
rect 124 275 126 277
rect 134 274 136 276
rect 134 267 136 269
rect 146 282 148 284
rect 146 275 148 277
rect 181 282 183 284
rect 169 263 171 265
rect 225 282 227 284
rect 225 275 227 277
rect 235 274 237 276
rect 235 267 237 269
rect 247 282 249 284
rect 247 275 249 277
rect 282 282 284 284
rect 270 263 272 265
rect 326 282 328 284
rect 326 275 328 277
rect 336 274 338 276
rect 336 267 338 269
rect 348 282 350 284
rect 348 275 350 277
rect 383 282 385 284
rect 371 263 373 265
rect 446 276 448 278
rect 479 282 481 284
rect 479 275 481 277
rect 489 274 491 276
rect 489 267 491 269
rect 501 282 503 284
rect 501 275 503 277
rect 536 282 538 284
rect 524 263 526 265
rect 580 282 582 284
rect 580 275 582 277
rect 590 274 592 276
rect 590 267 592 269
rect 602 282 604 284
rect 602 275 604 277
rect 637 282 639 284
rect 625 263 627 265
rect 679 282 681 284
rect 679 275 681 277
rect 689 274 691 276
rect 689 267 691 269
rect 701 282 703 284
rect 701 275 703 277
rect 736 282 738 284
rect 724 263 726 265
<< pdifct1 >>
rect 103 563 105 565
rect 103 556 105 558
rect 143 563 145 565
rect 143 556 145 558
rect 154 555 156 557
rect 154 548 156 550
rect 232 558 234 560
rect 232 551 234 553
rect 250 558 252 560
rect 250 551 252 553
rect 339 563 341 565
rect 328 555 330 557
rect 339 556 341 558
rect 328 548 330 550
rect 379 563 381 565
rect 379 556 381 558
rect 420 558 422 560
rect 420 551 422 553
rect 509 563 511 565
rect 498 555 500 557
rect 509 556 511 558
rect 498 548 500 550
rect 549 563 551 565
rect 549 556 551 558
rect 619 563 621 565
rect 619 556 621 558
rect 659 563 661 565
rect 659 556 661 558
rect 670 555 672 557
rect 670 548 672 550
rect 748 558 750 560
rect 748 551 750 553
rect 103 458 105 460
rect 103 451 105 453
rect 154 466 156 468
rect 143 458 145 460
rect 143 451 145 453
rect 232 463 234 465
rect 232 456 234 458
rect 250 463 252 465
rect 250 456 252 458
rect 328 466 330 468
rect 328 459 330 461
rect 339 458 341 460
rect 339 451 341 453
rect 379 458 381 460
rect 379 451 381 453
rect 420 463 422 465
rect 420 456 422 458
rect 498 466 500 468
rect 498 459 500 461
rect 509 458 511 460
rect 509 451 511 453
rect 549 458 551 460
rect 549 451 551 453
rect 619 458 621 460
rect 619 451 621 453
rect 670 466 672 468
rect 659 458 661 460
rect 670 459 672 461
rect 659 451 661 453
rect 748 463 750 465
rect 748 456 750 458
rect 73 420 75 422
rect 73 413 75 415
rect 84 429 86 431
rect 114 411 116 413
rect 114 404 116 406
rect 192 414 194 416
rect 192 407 194 409
rect 215 411 217 413
rect 215 404 217 406
rect 293 414 295 416
rect 293 407 295 409
rect 317 411 319 413
rect 317 404 319 406
rect 417 420 419 422
rect 395 414 397 416
rect 417 413 419 415
rect 395 407 397 409
rect 428 429 430 431
rect 470 411 472 413
rect 470 404 472 406
rect 548 414 550 416
rect 548 407 550 409
rect 571 411 573 413
rect 571 404 573 406
rect 649 414 651 416
rect 649 407 651 409
rect 670 411 672 413
rect 670 404 672 406
rect 748 414 750 416
rect 748 407 750 409
rect 75 322 77 324
rect 75 315 77 317
rect 153 319 155 321
rect 153 312 155 314
rect 163 313 165 315
rect 163 306 165 308
rect 174 297 176 299
rect 216 322 218 324
rect 216 315 218 317
rect 294 319 296 321
rect 294 312 296 314
rect 316 319 318 321
rect 316 312 318 314
rect 394 322 396 324
rect 394 315 396 317
rect 417 313 419 315
rect 417 306 419 308
rect 428 297 430 299
rect 470 322 472 324
rect 470 315 472 317
rect 548 319 550 321
rect 548 312 550 314
rect 571 322 573 324
rect 571 315 573 317
rect 649 319 651 321
rect 649 312 651 314
rect 670 322 672 324
rect 670 315 672 317
rect 748 319 750 321
rect 748 312 750 314
rect 73 276 75 278
rect 73 269 75 271
rect 84 285 86 287
rect 114 267 116 269
rect 114 260 116 262
rect 192 270 194 272
rect 192 263 194 265
rect 215 267 217 269
rect 215 260 217 262
rect 293 270 295 272
rect 293 263 295 265
rect 316 267 318 269
rect 316 260 318 262
rect 416 276 418 278
rect 394 270 396 272
rect 416 269 418 271
rect 394 263 396 265
rect 427 285 429 287
rect 469 267 471 269
rect 469 260 471 262
rect 547 270 549 272
rect 547 263 549 265
rect 570 267 572 269
rect 570 260 572 262
rect 648 270 650 272
rect 648 263 650 265
rect 669 267 671 269
rect 669 260 671 262
rect 747 270 749 272
rect 747 263 749 265
<< alu0 >>
rect 71 570 73 572
rect 75 570 77 572
rect 71 565 77 570
rect 91 570 93 572
rect 95 570 97 572
rect 71 563 73 565
rect 75 563 77 565
rect 71 562 77 563
rect 81 566 87 567
rect 81 564 83 566
rect 85 564 87 566
rect 81 559 87 564
rect 91 565 97 570
rect 111 570 113 572
rect 115 570 117 572
rect 91 563 93 565
rect 95 563 97 565
rect 91 562 97 563
rect 81 557 83 559
rect 85 558 87 559
rect 111 565 117 570
rect 131 570 133 572
rect 135 570 137 572
rect 111 563 113 565
rect 115 563 117 565
rect 111 562 117 563
rect 121 566 127 567
rect 121 564 123 566
rect 125 564 127 566
rect 121 559 127 564
rect 131 565 137 570
rect 162 570 164 572
rect 166 570 168 572
rect 131 563 133 565
rect 135 563 137 565
rect 131 562 137 563
rect 85 557 95 558
rect 81 554 95 557
rect 91 550 95 554
rect 91 546 99 550
rect 95 541 99 546
rect 95 539 96 541
rect 98 539 99 541
rect 95 534 99 539
rect 87 530 99 534
rect 87 526 91 530
rect 102 527 103 534
rect 121 557 123 559
rect 125 558 127 559
rect 162 565 168 570
rect 184 570 186 572
rect 188 570 190 572
rect 162 563 164 565
rect 166 563 168 565
rect 162 562 168 563
rect 173 564 177 566
rect 173 562 174 564
rect 176 562 177 564
rect 184 565 190 570
rect 219 570 221 572
rect 223 570 225 572
rect 219 569 225 570
rect 259 570 261 572
rect 263 570 265 572
rect 259 569 265 570
rect 294 570 296 572
rect 298 570 300 572
rect 184 563 186 565
rect 188 563 190 565
rect 184 562 190 563
rect 125 557 135 558
rect 121 554 135 557
rect 131 550 135 554
rect 131 546 139 550
rect 135 541 139 546
rect 135 539 136 541
rect 138 539 139 541
rect 135 534 139 539
rect 127 530 139 534
rect 71 525 91 526
rect 71 523 73 525
rect 75 523 91 525
rect 71 522 91 523
rect 127 526 131 530
rect 142 527 143 534
rect 111 525 131 526
rect 111 523 113 525
rect 115 523 131 525
rect 111 522 131 523
rect 173 558 177 562
rect 196 558 220 562
rect 160 557 200 558
rect 160 555 174 557
rect 176 555 200 557
rect 160 554 200 555
rect 160 543 164 554
rect 208 553 212 555
rect 216 554 222 558
rect 208 551 209 553
rect 211 551 212 553
rect 208 550 212 551
rect 208 546 215 550
rect 158 541 164 543
rect 158 539 159 541
rect 161 539 164 541
rect 158 537 164 539
rect 168 541 172 546
rect 168 539 169 541
rect 171 539 172 541
rect 168 537 172 539
rect 160 534 164 537
rect 160 530 180 534
rect 176 526 180 530
rect 211 535 215 546
rect 218 544 222 554
rect 218 542 219 544
rect 221 542 222 544
rect 218 540 222 542
rect 211 534 229 535
rect 191 532 195 534
rect 211 533 225 534
rect 191 530 192 532
rect 194 530 195 532
rect 176 525 186 526
rect 176 523 182 525
rect 184 523 186 525
rect 176 522 186 523
rect 191 525 195 530
rect 200 532 225 533
rect 227 532 229 534
rect 200 530 202 532
rect 204 531 229 532
rect 204 530 215 531
rect 200 529 215 530
rect 191 523 192 525
rect 194 524 216 525
rect 194 523 212 524
rect 191 522 212 523
rect 214 522 216 524
rect 191 521 216 522
rect 221 521 225 523
rect 294 565 300 570
rect 316 570 318 572
rect 320 570 322 572
rect 294 563 296 565
rect 298 563 300 565
rect 294 562 300 563
rect 307 564 311 566
rect 307 562 308 564
rect 310 562 311 564
rect 316 565 322 570
rect 347 570 349 572
rect 351 570 353 572
rect 316 563 318 565
rect 320 563 322 565
rect 316 562 322 563
rect 264 558 288 562
rect 307 558 311 562
rect 262 554 268 558
rect 284 557 324 558
rect 284 555 308 557
rect 310 555 324 557
rect 262 544 266 554
rect 272 553 276 555
rect 284 554 324 555
rect 272 551 273 553
rect 275 551 276 553
rect 272 550 276 551
rect 262 542 263 544
rect 265 542 266 544
rect 262 540 266 542
rect 269 546 276 550
rect 269 535 273 546
rect 312 541 316 546
rect 312 539 313 541
rect 315 539 316 541
rect 255 534 273 535
rect 255 532 257 534
rect 259 533 273 534
rect 259 532 284 533
rect 255 531 280 532
rect 269 530 280 531
rect 282 530 284 532
rect 269 529 284 530
rect 289 532 293 534
rect 289 530 290 532
rect 292 530 293 532
rect 289 525 293 530
rect 312 537 316 539
rect 320 543 324 554
rect 320 541 326 543
rect 320 539 323 541
rect 325 539 326 541
rect 320 537 326 539
rect 320 534 324 537
rect 304 530 324 534
rect 304 526 308 530
rect 268 524 290 525
rect 259 521 263 523
rect 268 522 270 524
rect 272 523 290 524
rect 292 523 293 525
rect 272 522 293 523
rect 298 525 308 526
rect 298 523 300 525
rect 302 523 308 525
rect 298 522 308 523
rect 347 565 353 570
rect 367 570 369 572
rect 371 570 373 572
rect 347 563 349 565
rect 351 563 353 565
rect 347 562 353 563
rect 357 566 363 567
rect 357 564 359 566
rect 361 564 363 566
rect 357 559 363 564
rect 367 565 373 570
rect 387 570 389 572
rect 391 570 393 572
rect 367 563 369 565
rect 371 563 373 565
rect 367 562 373 563
rect 357 558 359 559
rect 349 557 359 558
rect 361 557 363 559
rect 349 554 363 557
rect 349 550 353 554
rect 345 546 353 550
rect 387 565 393 570
rect 407 570 409 572
rect 411 570 413 572
rect 387 563 389 565
rect 391 563 393 565
rect 387 562 393 563
rect 397 566 403 567
rect 397 564 399 566
rect 401 564 403 566
rect 397 559 403 564
rect 407 565 413 570
rect 429 570 431 572
rect 433 570 435 572
rect 429 569 435 570
rect 464 570 466 572
rect 468 570 470 572
rect 407 563 409 565
rect 411 563 413 565
rect 407 562 413 563
rect 464 565 470 570
rect 486 570 488 572
rect 490 570 492 572
rect 464 563 466 565
rect 468 563 470 565
rect 464 562 470 563
rect 477 564 481 566
rect 477 562 478 564
rect 480 562 481 564
rect 486 565 492 570
rect 517 570 519 572
rect 521 570 523 572
rect 486 563 488 565
rect 490 563 492 565
rect 486 562 492 563
rect 397 558 399 559
rect 389 557 399 558
rect 401 557 403 559
rect 389 554 403 557
rect 345 541 349 546
rect 345 539 346 541
rect 348 539 349 541
rect 345 534 349 539
rect 341 527 342 534
rect 345 530 357 534
rect 353 526 357 530
rect 389 550 393 554
rect 385 546 393 550
rect 434 558 458 562
rect 477 558 481 562
rect 432 554 438 558
rect 454 557 494 558
rect 454 555 478 557
rect 480 555 494 557
rect 385 541 389 546
rect 385 539 386 541
rect 388 539 389 541
rect 385 534 389 539
rect 381 527 382 534
rect 385 530 397 534
rect 353 525 373 526
rect 353 523 369 525
rect 371 523 373 525
rect 353 522 373 523
rect 393 526 397 530
rect 432 544 436 554
rect 442 553 446 555
rect 454 554 494 555
rect 442 551 443 553
rect 445 551 446 553
rect 442 550 446 551
rect 432 542 433 544
rect 435 542 436 544
rect 432 540 436 542
rect 439 546 446 550
rect 439 535 443 546
rect 482 541 486 546
rect 482 539 483 541
rect 485 539 486 541
rect 425 534 443 535
rect 425 532 427 534
rect 429 533 443 534
rect 429 532 454 533
rect 425 531 450 532
rect 439 530 450 531
rect 452 530 454 532
rect 439 529 454 530
rect 459 532 463 534
rect 459 530 460 532
rect 462 530 463 532
rect 393 525 413 526
rect 393 523 409 525
rect 411 523 413 525
rect 393 522 413 523
rect 459 525 463 530
rect 482 537 486 539
rect 490 543 494 554
rect 490 541 496 543
rect 490 539 493 541
rect 495 539 496 541
rect 490 537 496 539
rect 490 534 494 537
rect 474 530 494 534
rect 474 526 478 530
rect 438 524 460 525
rect 268 521 293 522
rect 429 521 433 523
rect 438 522 440 524
rect 442 523 460 524
rect 462 523 463 525
rect 442 522 463 523
rect 468 525 478 526
rect 468 523 470 525
rect 472 523 478 525
rect 468 522 478 523
rect 517 565 523 570
rect 537 570 539 572
rect 541 570 543 572
rect 517 563 519 565
rect 521 563 523 565
rect 517 562 523 563
rect 527 566 533 567
rect 527 564 529 566
rect 531 564 533 566
rect 527 559 533 564
rect 537 565 543 570
rect 557 570 559 572
rect 561 570 563 572
rect 537 563 539 565
rect 541 563 543 565
rect 537 562 543 563
rect 527 558 529 559
rect 519 557 529 558
rect 531 557 533 559
rect 519 554 533 557
rect 519 550 523 554
rect 515 546 523 550
rect 557 565 563 570
rect 577 570 579 572
rect 581 570 583 572
rect 557 563 559 565
rect 561 563 563 565
rect 557 562 563 563
rect 567 566 573 567
rect 567 564 569 566
rect 571 564 573 566
rect 567 559 573 564
rect 577 565 583 570
rect 577 563 579 565
rect 581 563 583 565
rect 577 562 583 563
rect 587 570 589 572
rect 591 570 593 572
rect 587 565 593 570
rect 607 570 609 572
rect 611 570 613 572
rect 587 563 589 565
rect 591 563 593 565
rect 587 562 593 563
rect 597 566 603 567
rect 597 564 599 566
rect 601 564 603 566
rect 597 559 603 564
rect 607 565 613 570
rect 627 570 629 572
rect 631 570 633 572
rect 607 563 609 565
rect 611 563 613 565
rect 607 562 613 563
rect 567 558 569 559
rect 559 557 569 558
rect 571 557 573 559
rect 559 554 573 557
rect 515 541 519 546
rect 515 539 516 541
rect 518 539 519 541
rect 515 534 519 539
rect 511 527 512 534
rect 515 530 527 534
rect 523 526 527 530
rect 559 550 563 554
rect 555 546 563 550
rect 597 557 599 559
rect 601 558 603 559
rect 627 565 633 570
rect 647 570 649 572
rect 651 570 653 572
rect 627 563 629 565
rect 631 563 633 565
rect 627 562 633 563
rect 637 566 643 567
rect 637 564 639 566
rect 641 564 643 566
rect 637 559 643 564
rect 647 565 653 570
rect 678 570 680 572
rect 682 570 684 572
rect 647 563 649 565
rect 651 563 653 565
rect 647 562 653 563
rect 601 557 611 558
rect 597 554 611 557
rect 607 550 611 554
rect 607 546 615 550
rect 555 541 559 546
rect 555 539 556 541
rect 558 539 559 541
rect 555 534 559 539
rect 551 527 552 534
rect 555 530 567 534
rect 523 525 543 526
rect 523 523 539 525
rect 541 523 543 525
rect 523 522 543 523
rect 563 526 567 530
rect 611 541 615 546
rect 611 539 612 541
rect 614 539 615 541
rect 611 534 615 539
rect 603 530 615 534
rect 603 526 607 530
rect 618 527 619 534
rect 637 557 639 559
rect 641 558 643 559
rect 678 565 684 570
rect 700 570 702 572
rect 704 570 706 572
rect 678 563 680 565
rect 682 563 684 565
rect 678 562 684 563
rect 689 564 693 566
rect 689 562 690 564
rect 692 562 693 564
rect 700 565 706 570
rect 735 570 737 572
rect 739 570 741 572
rect 735 569 741 570
rect 700 563 702 565
rect 704 563 706 565
rect 700 562 706 563
rect 641 557 651 558
rect 637 554 651 557
rect 647 550 651 554
rect 647 546 655 550
rect 651 541 655 546
rect 651 539 652 541
rect 654 539 655 541
rect 651 534 655 539
rect 643 530 655 534
rect 563 525 583 526
rect 563 523 579 525
rect 581 523 583 525
rect 563 522 583 523
rect 587 525 607 526
rect 587 523 589 525
rect 591 523 607 525
rect 587 522 607 523
rect 643 526 647 530
rect 658 527 659 534
rect 627 525 647 526
rect 627 523 629 525
rect 631 523 647 525
rect 627 522 647 523
rect 689 558 693 562
rect 712 558 736 562
rect 676 557 716 558
rect 676 555 690 557
rect 692 555 716 557
rect 676 554 716 555
rect 676 543 680 554
rect 724 553 728 555
rect 732 554 738 558
rect 724 551 725 553
rect 727 551 728 553
rect 724 550 728 551
rect 724 546 731 550
rect 674 541 680 543
rect 674 539 675 541
rect 677 539 680 541
rect 674 537 680 539
rect 684 541 688 546
rect 684 539 685 541
rect 687 539 688 541
rect 684 537 688 539
rect 676 534 680 537
rect 676 530 696 534
rect 692 526 696 530
rect 727 535 731 546
rect 734 544 738 554
rect 734 542 735 544
rect 737 542 738 544
rect 734 540 738 542
rect 727 534 745 535
rect 707 532 711 534
rect 727 533 741 534
rect 707 530 708 532
rect 710 530 711 532
rect 692 525 702 526
rect 692 523 698 525
rect 700 523 702 525
rect 692 522 702 523
rect 707 525 711 530
rect 716 532 741 533
rect 743 532 745 534
rect 716 530 718 532
rect 720 531 745 532
rect 720 530 731 531
rect 716 529 731 530
rect 707 523 708 525
rect 710 524 732 525
rect 710 523 728 524
rect 707 522 728 523
rect 730 522 732 524
rect 438 521 463 522
rect 707 521 732 522
rect 737 521 741 523
rect 221 519 222 521
rect 224 519 225 521
rect 163 518 169 519
rect 163 516 165 518
rect 167 516 169 518
rect 221 516 225 519
rect 259 519 260 521
rect 262 519 263 521
rect 429 519 430 521
rect 432 519 433 521
rect 737 519 738 521
rect 740 519 741 521
rect 259 516 263 519
rect 315 518 321 519
rect 315 516 317 518
rect 319 516 321 518
rect 429 516 433 519
rect 485 518 491 519
rect 485 516 487 518
rect 489 516 491 518
rect 679 518 685 519
rect 679 516 681 518
rect 683 516 685 518
rect 737 516 741 519
rect 163 498 165 500
rect 167 498 169 500
rect 163 497 169 498
rect 221 497 225 500
rect 221 495 222 497
rect 224 495 225 497
rect 259 497 263 500
rect 315 498 317 500
rect 319 498 321 500
rect 315 497 321 498
rect 429 497 433 500
rect 485 498 487 500
rect 489 498 491 500
rect 485 497 491 498
rect 679 498 681 500
rect 683 498 685 500
rect 679 497 685 498
rect 737 497 741 500
rect 259 495 260 497
rect 262 495 263 497
rect 429 495 430 497
rect 432 495 433 497
rect 737 495 738 497
rect 740 495 741 497
rect 191 494 216 495
rect 71 493 91 494
rect 71 491 73 493
rect 75 491 91 493
rect 71 490 91 491
rect 87 486 91 490
rect 111 493 131 494
rect 111 491 113 493
rect 115 491 131 493
rect 111 490 131 491
rect 87 482 99 486
rect 102 482 103 489
rect 95 477 99 482
rect 95 475 96 477
rect 98 475 99 477
rect 95 470 99 475
rect 91 466 99 470
rect 91 462 95 466
rect 127 486 131 490
rect 127 482 139 486
rect 142 482 143 489
rect 135 477 139 482
rect 135 475 136 477
rect 138 475 139 477
rect 135 470 139 475
rect 81 459 95 462
rect 81 457 83 459
rect 85 458 95 459
rect 85 457 87 458
rect 71 453 77 454
rect 71 451 73 453
rect 75 451 77 453
rect 71 446 77 451
rect 81 452 87 457
rect 81 450 83 452
rect 85 450 87 452
rect 81 449 87 450
rect 91 453 97 454
rect 91 451 93 453
rect 95 451 97 453
rect 71 444 73 446
rect 75 444 77 446
rect 91 446 97 451
rect 131 466 139 470
rect 131 462 135 466
rect 121 459 135 462
rect 121 457 123 459
rect 125 458 135 459
rect 125 457 127 458
rect 111 453 117 454
rect 111 451 113 453
rect 115 451 117 453
rect 91 444 93 446
rect 95 444 97 446
rect 111 446 117 451
rect 121 452 127 457
rect 121 450 123 452
rect 125 450 127 452
rect 121 449 127 450
rect 131 453 137 454
rect 131 451 133 453
rect 135 451 137 453
rect 111 444 113 446
rect 115 444 117 446
rect 131 446 137 451
rect 176 493 186 494
rect 176 491 182 493
rect 184 491 186 493
rect 176 490 186 491
rect 191 493 212 494
rect 191 491 192 493
rect 194 492 212 493
rect 214 492 216 494
rect 221 493 225 495
rect 194 491 216 492
rect 176 486 180 490
rect 160 482 180 486
rect 160 479 164 482
rect 158 477 164 479
rect 158 475 159 477
rect 161 475 164 477
rect 158 473 164 475
rect 160 462 164 473
rect 168 477 172 479
rect 191 486 195 491
rect 191 484 192 486
rect 194 484 195 486
rect 191 482 195 484
rect 200 486 215 487
rect 200 484 202 486
rect 204 485 215 486
rect 204 484 229 485
rect 200 483 225 484
rect 211 482 225 483
rect 227 482 229 484
rect 211 481 229 482
rect 168 475 169 477
rect 171 475 172 477
rect 168 470 172 475
rect 211 470 215 481
rect 208 466 215 470
rect 218 474 222 476
rect 218 472 219 474
rect 221 472 222 474
rect 208 465 212 466
rect 208 463 209 465
rect 211 463 212 465
rect 160 461 200 462
rect 208 461 212 463
rect 218 462 222 472
rect 160 459 174 461
rect 176 459 200 461
rect 160 458 200 459
rect 216 458 222 462
rect 173 454 177 458
rect 196 454 220 458
rect 162 453 168 454
rect 162 451 164 453
rect 166 451 168 453
rect 131 444 133 446
rect 135 444 137 446
rect 162 446 168 451
rect 173 452 174 454
rect 176 452 177 454
rect 173 450 177 452
rect 184 453 190 454
rect 184 451 186 453
rect 188 451 190 453
rect 162 444 164 446
rect 166 444 168 446
rect 184 446 190 451
rect 259 493 263 495
rect 268 494 293 495
rect 268 492 270 494
rect 272 493 293 494
rect 272 492 290 493
rect 268 491 290 492
rect 292 491 293 493
rect 269 486 284 487
rect 269 485 280 486
rect 255 484 280 485
rect 282 484 284 486
rect 255 482 257 484
rect 259 483 284 484
rect 289 486 293 491
rect 298 493 308 494
rect 298 491 300 493
rect 302 491 308 493
rect 298 490 308 491
rect 289 484 290 486
rect 292 484 293 486
rect 259 482 273 483
rect 289 482 293 484
rect 255 481 273 482
rect 262 474 266 476
rect 262 472 263 474
rect 265 472 266 474
rect 262 462 266 472
rect 269 470 273 481
rect 304 486 308 490
rect 304 482 324 486
rect 320 479 324 482
rect 312 477 316 479
rect 312 475 313 477
rect 315 475 316 477
rect 312 470 316 475
rect 320 477 326 479
rect 320 475 323 477
rect 325 475 326 477
rect 320 473 326 475
rect 269 466 276 470
rect 272 465 276 466
rect 272 463 273 465
rect 275 463 276 465
rect 262 458 268 462
rect 272 461 276 463
rect 320 462 324 473
rect 284 461 324 462
rect 284 459 308 461
rect 310 459 324 461
rect 284 458 324 459
rect 264 454 288 458
rect 307 454 311 458
rect 353 493 373 494
rect 353 491 369 493
rect 371 491 373 493
rect 353 490 373 491
rect 341 482 342 489
rect 353 486 357 490
rect 393 493 413 494
rect 393 491 409 493
rect 411 491 413 493
rect 393 490 413 491
rect 429 493 433 495
rect 438 494 463 495
rect 707 494 732 495
rect 438 492 440 494
rect 442 493 463 494
rect 442 492 460 493
rect 438 491 460 492
rect 462 491 463 493
rect 345 482 357 486
rect 345 477 349 482
rect 345 475 346 477
rect 348 475 349 477
rect 345 470 349 475
rect 345 466 353 470
rect 349 462 353 466
rect 349 459 363 462
rect 349 458 359 459
rect 294 453 300 454
rect 294 451 296 453
rect 298 451 300 453
rect 184 444 186 446
rect 188 444 190 446
rect 219 446 225 447
rect 219 444 221 446
rect 223 444 225 446
rect 259 446 265 447
rect 259 444 261 446
rect 263 444 265 446
rect 294 446 300 451
rect 307 452 308 454
rect 310 452 311 454
rect 307 450 311 452
rect 316 453 322 454
rect 316 451 318 453
rect 320 451 322 453
rect 294 444 296 446
rect 298 444 300 446
rect 316 446 322 451
rect 357 457 359 458
rect 361 457 363 459
rect 381 482 382 489
rect 393 486 397 490
rect 385 482 397 486
rect 385 477 389 482
rect 385 475 386 477
rect 388 475 389 477
rect 385 470 389 475
rect 385 466 393 470
rect 389 462 393 466
rect 389 459 403 462
rect 389 458 399 459
rect 347 453 353 454
rect 347 451 349 453
rect 351 451 353 453
rect 316 444 318 446
rect 320 444 322 446
rect 347 446 353 451
rect 357 452 363 457
rect 397 457 399 458
rect 401 457 403 459
rect 439 486 454 487
rect 439 485 450 486
rect 425 484 450 485
rect 452 484 454 486
rect 425 482 427 484
rect 429 483 454 484
rect 459 486 463 491
rect 468 493 478 494
rect 468 491 470 493
rect 472 491 478 493
rect 468 490 478 491
rect 459 484 460 486
rect 462 484 463 486
rect 429 482 443 483
rect 459 482 463 484
rect 425 481 443 482
rect 432 474 436 476
rect 432 472 433 474
rect 435 472 436 474
rect 432 462 436 472
rect 439 470 443 481
rect 474 486 478 490
rect 474 482 494 486
rect 490 479 494 482
rect 482 477 486 479
rect 482 475 483 477
rect 485 475 486 477
rect 482 470 486 475
rect 490 477 496 479
rect 490 475 493 477
rect 495 475 496 477
rect 490 473 496 475
rect 439 466 446 470
rect 442 465 446 466
rect 442 463 443 465
rect 445 463 446 465
rect 432 458 438 462
rect 442 461 446 463
rect 490 462 494 473
rect 454 461 494 462
rect 454 459 478 461
rect 480 459 494 461
rect 454 458 494 459
rect 357 450 359 452
rect 361 450 363 452
rect 357 449 363 450
rect 367 453 373 454
rect 367 451 369 453
rect 371 451 373 453
rect 347 444 349 446
rect 351 444 353 446
rect 367 446 373 451
rect 387 453 393 454
rect 387 451 389 453
rect 391 451 393 453
rect 367 444 369 446
rect 371 444 373 446
rect 387 446 393 451
rect 397 452 403 457
rect 434 454 458 458
rect 477 454 481 458
rect 523 493 543 494
rect 523 491 539 493
rect 541 491 543 493
rect 523 490 543 491
rect 511 482 512 489
rect 523 486 527 490
rect 563 493 583 494
rect 563 491 579 493
rect 581 491 583 493
rect 563 490 583 491
rect 587 493 607 494
rect 587 491 589 493
rect 591 491 607 493
rect 587 490 607 491
rect 515 482 527 486
rect 515 477 519 482
rect 515 475 516 477
rect 518 475 519 477
rect 515 470 519 475
rect 551 482 552 489
rect 563 486 567 490
rect 555 482 567 486
rect 515 466 523 470
rect 519 462 523 466
rect 519 459 533 462
rect 519 458 529 459
rect 397 450 399 452
rect 401 450 403 452
rect 397 449 403 450
rect 407 453 413 454
rect 407 451 409 453
rect 411 451 413 453
rect 387 444 389 446
rect 391 444 393 446
rect 407 446 413 451
rect 464 453 470 454
rect 464 451 466 453
rect 468 451 470 453
rect 407 444 409 446
rect 411 444 413 446
rect 429 446 435 447
rect 429 444 431 446
rect 433 444 435 446
rect 464 446 470 451
rect 477 452 478 454
rect 480 452 481 454
rect 477 450 481 452
rect 486 453 492 454
rect 486 451 488 453
rect 490 451 492 453
rect 464 444 466 446
rect 468 444 470 446
rect 486 446 492 451
rect 527 457 529 458
rect 531 457 533 459
rect 555 477 559 482
rect 555 475 556 477
rect 558 475 559 477
rect 555 470 559 475
rect 603 486 607 490
rect 627 493 647 494
rect 627 491 629 493
rect 631 491 647 493
rect 627 490 647 491
rect 603 482 615 486
rect 618 482 619 489
rect 611 477 615 482
rect 611 475 612 477
rect 614 475 615 477
rect 611 470 615 475
rect 555 466 563 470
rect 559 462 563 466
rect 559 459 573 462
rect 559 458 569 459
rect 517 453 523 454
rect 517 451 519 453
rect 521 451 523 453
rect 486 444 488 446
rect 490 444 492 446
rect 517 446 523 451
rect 527 452 533 457
rect 527 450 529 452
rect 531 450 533 452
rect 527 449 533 450
rect 537 453 543 454
rect 537 451 539 453
rect 541 451 543 453
rect 517 444 519 446
rect 521 444 523 446
rect 537 446 543 451
rect 567 457 569 458
rect 571 457 573 459
rect 607 466 615 470
rect 607 462 611 466
rect 643 486 647 490
rect 643 482 655 486
rect 658 482 659 489
rect 651 477 655 482
rect 651 475 652 477
rect 654 475 655 477
rect 651 470 655 475
rect 597 459 611 462
rect 597 457 599 459
rect 601 458 611 459
rect 601 457 603 458
rect 557 453 563 454
rect 557 451 559 453
rect 561 451 563 453
rect 537 444 539 446
rect 541 444 543 446
rect 557 446 563 451
rect 567 452 573 457
rect 567 450 569 452
rect 571 450 573 452
rect 567 449 573 450
rect 577 453 583 454
rect 577 451 579 453
rect 581 451 583 453
rect 557 444 559 446
rect 561 444 563 446
rect 577 446 583 451
rect 577 444 579 446
rect 581 444 583 446
rect 587 453 593 454
rect 587 451 589 453
rect 591 451 593 453
rect 587 446 593 451
rect 597 452 603 457
rect 597 450 599 452
rect 601 450 603 452
rect 597 449 603 450
rect 607 453 613 454
rect 607 451 609 453
rect 611 451 613 453
rect 587 444 589 446
rect 591 444 593 446
rect 607 446 613 451
rect 647 466 655 470
rect 647 462 651 466
rect 637 459 651 462
rect 637 457 639 459
rect 641 458 651 459
rect 641 457 643 458
rect 627 453 633 454
rect 627 451 629 453
rect 631 451 633 453
rect 607 444 609 446
rect 611 444 613 446
rect 627 446 633 451
rect 637 452 643 457
rect 637 450 639 452
rect 641 450 643 452
rect 637 449 643 450
rect 647 453 653 454
rect 647 451 649 453
rect 651 451 653 453
rect 627 444 629 446
rect 631 444 633 446
rect 647 446 653 451
rect 692 493 702 494
rect 692 491 698 493
rect 700 491 702 493
rect 692 490 702 491
rect 707 493 728 494
rect 707 491 708 493
rect 710 492 728 493
rect 730 492 732 494
rect 737 493 741 495
rect 710 491 732 492
rect 692 486 696 490
rect 676 482 696 486
rect 676 479 680 482
rect 674 477 680 479
rect 674 475 675 477
rect 677 475 680 477
rect 674 473 680 475
rect 676 462 680 473
rect 684 477 688 479
rect 707 486 711 491
rect 707 484 708 486
rect 710 484 711 486
rect 707 482 711 484
rect 716 486 731 487
rect 716 484 718 486
rect 720 485 731 486
rect 720 484 745 485
rect 716 483 741 484
rect 727 482 741 483
rect 743 482 745 484
rect 727 481 745 482
rect 684 475 685 477
rect 687 475 688 477
rect 684 470 688 475
rect 727 470 731 481
rect 724 466 731 470
rect 734 474 738 476
rect 734 472 735 474
rect 737 472 738 474
rect 724 465 728 466
rect 724 463 725 465
rect 727 463 728 465
rect 676 461 716 462
rect 724 461 728 463
rect 734 462 738 472
rect 676 459 690 461
rect 692 459 716 461
rect 676 458 716 459
rect 732 458 738 462
rect 689 454 693 458
rect 712 454 736 458
rect 678 453 684 454
rect 678 451 680 453
rect 682 451 684 453
rect 647 444 649 446
rect 651 444 653 446
rect 678 446 684 451
rect 689 452 690 454
rect 692 452 693 454
rect 689 450 693 452
rect 700 453 706 454
rect 700 451 702 453
rect 704 451 706 453
rect 678 444 680 446
rect 682 444 684 446
rect 700 446 706 451
rect 700 444 702 446
rect 704 444 706 446
rect 735 446 741 447
rect 735 444 737 446
rect 739 444 741 446
rect 122 426 124 428
rect 126 426 128 428
rect 87 422 107 423
rect 87 420 103 422
rect 105 420 107 422
rect 87 419 107 420
rect 122 421 128 426
rect 144 426 146 428
rect 148 426 150 428
rect 122 419 124 421
rect 126 419 128 421
rect 75 411 76 417
rect 87 414 91 419
rect 122 418 128 419
rect 133 420 137 422
rect 133 418 134 420
rect 136 418 137 420
rect 144 421 150 426
rect 179 426 181 428
rect 183 426 185 428
rect 179 425 185 426
rect 223 426 225 428
rect 227 426 229 428
rect 144 419 146 421
rect 148 419 150 421
rect 144 418 150 419
rect 223 421 229 426
rect 245 426 247 428
rect 249 426 251 428
rect 223 419 225 421
rect 227 419 229 421
rect 223 418 229 419
rect 234 420 238 422
rect 234 418 235 420
rect 237 418 238 420
rect 245 421 251 426
rect 280 426 282 428
rect 284 426 286 428
rect 280 425 286 426
rect 325 426 327 428
rect 329 426 331 428
rect 245 419 247 421
rect 249 419 251 421
rect 245 418 251 419
rect 325 421 331 426
rect 347 426 349 428
rect 351 426 353 428
rect 325 419 327 421
rect 329 419 331 421
rect 325 418 331 419
rect 336 420 340 422
rect 336 418 337 420
rect 339 418 340 420
rect 347 421 353 426
rect 382 426 384 428
rect 386 426 388 428
rect 382 425 388 426
rect 478 426 480 428
rect 482 426 484 428
rect 347 419 349 421
rect 351 419 353 421
rect 347 418 353 419
rect 79 410 91 414
rect 133 414 137 418
rect 156 414 180 418
rect 79 397 83 410
rect 79 395 80 397
rect 82 395 83 397
rect 79 389 83 395
rect 102 393 103 409
rect 120 413 160 414
rect 120 411 134 413
rect 136 411 160 413
rect 120 410 160 411
rect 79 385 96 389
rect 92 383 96 385
rect 81 381 87 382
rect 81 379 83 381
rect 85 379 87 381
rect 92 381 93 383
rect 95 381 96 383
rect 92 379 96 381
rect 101 383 107 384
rect 101 381 103 383
rect 105 381 107 383
rect 81 372 87 379
rect 101 372 107 381
rect 120 399 124 410
rect 168 409 172 411
rect 176 410 182 414
rect 168 407 169 409
rect 171 407 172 409
rect 168 406 172 407
rect 168 402 175 406
rect 118 397 124 399
rect 118 395 119 397
rect 121 395 124 397
rect 118 393 124 395
rect 128 397 132 402
rect 128 395 129 397
rect 131 395 132 397
rect 128 393 132 395
rect 120 390 124 393
rect 120 386 140 390
rect 136 382 140 386
rect 171 391 175 402
rect 178 400 182 410
rect 178 398 179 400
rect 181 398 182 400
rect 178 396 182 398
rect 171 390 189 391
rect 151 388 155 390
rect 171 389 185 390
rect 151 386 152 388
rect 154 386 155 388
rect 136 381 146 382
rect 136 379 142 381
rect 144 379 146 381
rect 136 378 146 379
rect 151 381 155 386
rect 160 388 185 389
rect 187 388 189 390
rect 160 386 162 388
rect 164 387 189 388
rect 164 386 175 387
rect 160 385 175 386
rect 151 379 152 381
rect 154 380 176 381
rect 154 379 172 380
rect 151 378 172 379
rect 174 378 176 380
rect 151 377 176 378
rect 181 377 185 379
rect 234 414 238 418
rect 257 414 281 418
rect 221 413 261 414
rect 221 411 235 413
rect 237 411 261 413
rect 221 410 261 411
rect 221 399 225 410
rect 269 409 273 411
rect 277 410 283 414
rect 269 407 270 409
rect 272 407 273 409
rect 269 406 273 407
rect 269 402 276 406
rect 219 397 225 399
rect 219 395 220 397
rect 222 395 225 397
rect 219 393 225 395
rect 229 397 233 402
rect 229 395 230 397
rect 232 395 233 397
rect 229 393 233 395
rect 221 390 225 393
rect 221 386 241 390
rect 237 382 241 386
rect 272 391 276 402
rect 279 400 283 410
rect 279 398 280 400
rect 282 398 283 400
rect 279 396 283 398
rect 272 390 290 391
rect 252 388 256 390
rect 272 389 286 390
rect 252 386 253 388
rect 255 386 256 388
rect 237 381 247 382
rect 237 379 243 381
rect 245 379 247 381
rect 237 378 247 379
rect 252 381 256 386
rect 261 388 286 389
rect 288 388 290 390
rect 261 386 263 388
rect 265 387 290 388
rect 265 386 276 387
rect 261 385 276 386
rect 252 379 253 381
rect 255 380 277 381
rect 255 379 273 380
rect 252 378 273 379
rect 275 378 277 380
rect 252 377 277 378
rect 282 377 286 379
rect 336 414 340 418
rect 359 414 383 418
rect 323 413 363 414
rect 323 411 337 413
rect 339 411 363 413
rect 323 410 363 411
rect 323 399 327 410
rect 371 409 375 411
rect 379 410 385 414
rect 371 407 372 409
rect 374 407 375 409
rect 371 406 375 407
rect 371 402 378 406
rect 321 397 327 399
rect 321 395 322 397
rect 324 395 327 397
rect 321 393 327 395
rect 331 397 335 402
rect 331 395 332 397
rect 334 395 335 397
rect 331 393 335 395
rect 323 390 327 393
rect 323 386 343 390
rect 339 382 343 386
rect 374 391 378 402
rect 381 400 385 410
rect 381 398 382 400
rect 384 398 385 400
rect 381 396 385 398
rect 374 390 392 391
rect 354 388 358 390
rect 374 389 388 390
rect 354 386 355 388
rect 357 386 358 388
rect 339 381 349 382
rect 339 379 345 381
rect 347 379 349 381
rect 339 378 349 379
rect 354 381 358 386
rect 363 388 388 389
rect 390 388 392 390
rect 363 386 365 388
rect 367 387 392 388
rect 367 386 378 387
rect 363 385 378 386
rect 354 379 355 381
rect 357 380 379 381
rect 357 379 375 380
rect 354 378 375 379
rect 377 378 379 380
rect 354 377 379 378
rect 384 377 388 379
rect 431 422 451 423
rect 431 420 447 422
rect 449 420 451 422
rect 431 419 451 420
rect 478 421 484 426
rect 500 426 502 428
rect 504 426 506 428
rect 478 419 480 421
rect 482 419 484 421
rect 419 411 420 417
rect 431 414 435 419
rect 478 418 484 419
rect 489 420 493 422
rect 489 418 490 420
rect 492 418 493 420
rect 500 421 506 426
rect 535 426 537 428
rect 539 426 541 428
rect 535 425 541 426
rect 579 426 581 428
rect 583 426 585 428
rect 500 419 502 421
rect 504 419 506 421
rect 500 418 506 419
rect 579 421 585 426
rect 601 426 603 428
rect 605 426 607 428
rect 579 419 581 421
rect 583 419 585 421
rect 579 418 585 419
rect 590 420 594 422
rect 590 418 591 420
rect 593 418 594 420
rect 601 421 607 426
rect 636 426 638 428
rect 640 426 642 428
rect 636 425 642 426
rect 678 426 680 428
rect 682 426 684 428
rect 601 419 603 421
rect 605 419 607 421
rect 601 418 607 419
rect 678 421 684 426
rect 700 426 702 428
rect 704 426 706 428
rect 678 419 680 421
rect 682 419 684 421
rect 678 418 684 419
rect 689 420 693 422
rect 689 418 690 420
rect 692 418 693 420
rect 700 421 706 426
rect 735 426 737 428
rect 739 426 741 428
rect 735 425 741 426
rect 700 419 702 421
rect 704 419 706 421
rect 700 418 706 419
rect 423 410 435 414
rect 489 414 493 418
rect 512 414 536 418
rect 423 397 427 410
rect 423 395 424 397
rect 426 395 427 397
rect 423 389 427 395
rect 446 393 447 409
rect 476 413 516 414
rect 476 411 490 413
rect 492 411 516 413
rect 476 410 516 411
rect 423 385 440 389
rect 436 383 440 385
rect 425 381 431 382
rect 425 379 427 381
rect 429 379 431 381
rect 436 381 437 383
rect 439 381 440 383
rect 436 379 440 381
rect 445 383 451 384
rect 445 381 447 383
rect 449 381 451 383
rect 181 375 182 377
rect 184 375 185 377
rect 282 375 283 377
rect 285 375 286 377
rect 384 375 385 377
rect 387 375 388 377
rect 123 374 129 375
rect 123 372 125 374
rect 127 372 129 374
rect 181 372 185 375
rect 224 374 230 375
rect 224 372 226 374
rect 228 372 230 374
rect 282 372 286 375
rect 326 374 332 375
rect 326 372 328 374
rect 330 372 332 374
rect 384 372 388 375
rect 425 372 431 379
rect 445 372 451 381
rect 476 399 480 410
rect 524 409 528 411
rect 532 410 538 414
rect 524 407 525 409
rect 527 407 528 409
rect 524 406 528 407
rect 524 402 531 406
rect 474 397 480 399
rect 474 395 475 397
rect 477 395 480 397
rect 474 393 480 395
rect 484 397 488 402
rect 484 395 485 397
rect 487 395 488 397
rect 484 393 488 395
rect 476 390 480 393
rect 476 386 496 390
rect 492 382 496 386
rect 527 391 531 402
rect 534 400 538 410
rect 534 398 535 400
rect 537 398 538 400
rect 534 396 538 398
rect 527 390 545 391
rect 507 388 511 390
rect 527 389 541 390
rect 507 386 508 388
rect 510 386 511 388
rect 492 381 502 382
rect 492 379 498 381
rect 500 379 502 381
rect 492 378 502 379
rect 507 381 511 386
rect 516 388 541 389
rect 543 388 545 390
rect 516 386 518 388
rect 520 387 545 388
rect 520 386 531 387
rect 516 385 531 386
rect 507 379 508 381
rect 510 380 532 381
rect 510 379 528 380
rect 507 378 528 379
rect 530 378 532 380
rect 507 377 532 378
rect 537 377 541 379
rect 590 414 594 418
rect 613 414 637 418
rect 577 413 617 414
rect 577 411 591 413
rect 593 411 617 413
rect 577 410 617 411
rect 577 399 581 410
rect 625 409 629 411
rect 633 410 639 414
rect 625 407 626 409
rect 628 407 629 409
rect 625 406 629 407
rect 625 402 632 406
rect 575 397 581 399
rect 575 395 576 397
rect 578 395 581 397
rect 575 393 581 395
rect 585 397 589 402
rect 585 395 586 397
rect 588 395 589 397
rect 585 393 589 395
rect 577 390 581 393
rect 577 386 597 390
rect 593 382 597 386
rect 628 391 632 402
rect 635 400 639 410
rect 635 398 636 400
rect 638 398 639 400
rect 635 396 639 398
rect 628 390 646 391
rect 608 388 612 390
rect 628 389 642 390
rect 608 386 609 388
rect 611 386 612 388
rect 593 381 603 382
rect 593 379 599 381
rect 601 379 603 381
rect 593 378 603 379
rect 608 381 612 386
rect 617 388 642 389
rect 644 388 646 390
rect 617 386 619 388
rect 621 387 646 388
rect 621 386 632 387
rect 617 385 632 386
rect 608 379 609 381
rect 611 380 633 381
rect 611 379 629 380
rect 608 378 629 379
rect 631 378 633 380
rect 608 377 633 378
rect 638 377 642 379
rect 689 414 693 418
rect 712 414 736 418
rect 676 413 716 414
rect 676 411 690 413
rect 692 411 716 413
rect 676 410 716 411
rect 676 399 680 410
rect 724 409 728 411
rect 732 410 738 414
rect 724 407 725 409
rect 727 407 728 409
rect 724 406 728 407
rect 724 402 731 406
rect 674 397 680 399
rect 674 395 675 397
rect 677 395 680 397
rect 674 393 680 395
rect 684 397 688 402
rect 684 395 685 397
rect 687 395 688 397
rect 684 393 688 395
rect 676 390 680 393
rect 676 386 696 390
rect 692 382 696 386
rect 727 391 731 402
rect 734 400 738 410
rect 734 398 735 400
rect 737 398 738 400
rect 734 396 738 398
rect 727 390 745 391
rect 707 388 711 390
rect 727 389 741 390
rect 707 386 708 388
rect 710 386 711 388
rect 692 381 702 382
rect 692 379 698 381
rect 700 379 702 381
rect 692 378 702 379
rect 707 381 711 386
rect 716 388 741 389
rect 743 388 745 390
rect 716 386 718 388
rect 720 387 745 388
rect 720 386 731 387
rect 716 385 731 386
rect 707 379 708 381
rect 710 380 732 381
rect 710 379 728 380
rect 707 378 728 379
rect 730 378 732 380
rect 707 377 732 378
rect 737 377 741 379
rect 537 375 538 377
rect 540 375 541 377
rect 638 375 639 377
rect 641 375 642 377
rect 737 375 738 377
rect 740 375 741 377
rect 479 374 485 375
rect 479 372 481 374
rect 483 372 485 374
rect 537 372 541 375
rect 580 374 586 375
rect 580 372 582 374
rect 584 372 586 374
rect 638 372 642 375
rect 679 374 685 375
rect 679 372 681 374
rect 683 372 685 374
rect 737 372 741 375
rect 84 354 86 356
rect 88 354 90 356
rect 84 353 90 354
rect 142 353 146 356
rect 142 351 143 353
rect 145 351 146 353
rect 112 350 137 351
rect 97 349 107 350
rect 97 347 103 349
rect 105 347 107 349
rect 97 346 107 347
rect 112 349 133 350
rect 112 347 113 349
rect 115 348 133 349
rect 135 348 137 350
rect 142 349 146 351
rect 115 347 137 348
rect 97 342 101 346
rect 81 338 101 342
rect 81 335 85 338
rect 79 333 85 335
rect 79 331 80 333
rect 82 331 85 333
rect 79 329 85 331
rect 81 318 85 329
rect 89 333 93 335
rect 112 342 116 347
rect 112 340 113 342
rect 115 340 116 342
rect 112 338 116 340
rect 121 342 136 343
rect 121 340 123 342
rect 125 341 136 342
rect 125 340 150 341
rect 121 339 146 340
rect 132 338 146 339
rect 148 338 150 340
rect 132 337 150 338
rect 89 331 90 333
rect 92 331 93 333
rect 89 326 93 331
rect 132 326 136 337
rect 129 322 136 326
rect 139 330 143 332
rect 139 328 140 330
rect 142 328 143 330
rect 129 321 133 322
rect 129 319 130 321
rect 132 319 133 321
rect 81 317 121 318
rect 129 317 133 319
rect 139 318 143 328
rect 81 315 95 317
rect 97 315 121 317
rect 81 314 121 315
rect 137 314 143 318
rect 94 310 98 314
rect 117 310 141 314
rect 83 309 89 310
rect 83 307 85 309
rect 87 307 89 309
rect 83 302 89 307
rect 94 308 95 310
rect 97 308 98 310
rect 94 306 98 308
rect 105 309 111 310
rect 105 307 107 309
rect 109 307 111 309
rect 83 300 85 302
rect 87 300 89 302
rect 105 302 111 307
rect 171 349 177 356
rect 171 347 173 349
rect 175 347 177 349
rect 171 346 177 347
rect 182 347 186 349
rect 182 345 183 347
rect 185 345 186 347
rect 182 343 186 345
rect 191 347 197 356
rect 225 354 227 356
rect 229 354 231 356
rect 225 353 231 354
rect 283 353 287 356
rect 283 351 284 353
rect 286 351 287 353
rect 325 353 329 356
rect 381 354 383 356
rect 385 354 387 356
rect 381 353 387 354
rect 325 351 326 353
rect 328 351 329 353
rect 253 350 278 351
rect 191 345 193 347
rect 195 345 197 347
rect 191 344 197 345
rect 238 349 248 350
rect 238 347 244 349
rect 246 347 248 349
rect 238 346 248 347
rect 253 349 274 350
rect 253 347 254 349
rect 256 348 274 349
rect 276 348 278 350
rect 283 349 287 351
rect 256 347 278 348
rect 169 339 186 343
rect 169 333 173 339
rect 238 342 242 346
rect 222 338 242 342
rect 222 335 226 338
rect 169 331 170 333
rect 172 331 173 333
rect 169 318 173 331
rect 192 319 193 335
rect 165 311 166 317
rect 169 314 181 318
rect 177 309 181 314
rect 220 333 226 335
rect 220 331 221 333
rect 223 331 226 333
rect 220 329 226 331
rect 222 318 226 329
rect 230 333 234 335
rect 253 342 257 347
rect 253 340 254 342
rect 256 340 257 342
rect 253 338 257 340
rect 262 342 277 343
rect 262 340 264 342
rect 266 341 277 342
rect 266 340 291 341
rect 262 339 287 340
rect 273 338 287 339
rect 289 338 291 340
rect 273 337 291 338
rect 230 331 231 333
rect 233 331 234 333
rect 230 326 234 331
rect 273 326 277 337
rect 270 322 277 326
rect 280 330 284 332
rect 280 328 281 330
rect 283 328 284 330
rect 270 321 274 322
rect 270 319 271 321
rect 273 319 274 321
rect 222 317 262 318
rect 270 317 274 319
rect 280 318 284 328
rect 222 315 236 317
rect 238 315 262 317
rect 222 314 262 315
rect 278 314 284 318
rect 235 310 239 314
rect 258 310 282 314
rect 224 309 230 310
rect 177 308 197 309
rect 177 306 193 308
rect 195 306 197 308
rect 177 305 197 306
rect 224 307 226 309
rect 228 307 230 309
rect 105 300 107 302
rect 109 300 111 302
rect 140 302 146 303
rect 140 300 142 302
rect 144 300 146 302
rect 224 302 230 307
rect 235 308 236 310
rect 238 308 239 310
rect 235 306 239 308
rect 246 309 252 310
rect 246 307 248 309
rect 250 307 252 309
rect 224 300 226 302
rect 228 300 230 302
rect 246 302 252 307
rect 325 349 329 351
rect 334 350 359 351
rect 334 348 336 350
rect 338 349 359 350
rect 338 348 356 349
rect 334 347 356 348
rect 358 347 359 349
rect 335 342 350 343
rect 335 341 346 342
rect 321 340 346 341
rect 348 340 350 342
rect 321 338 323 340
rect 325 339 350 340
rect 355 342 359 347
rect 364 349 374 350
rect 364 347 366 349
rect 368 347 374 349
rect 364 346 374 347
rect 355 340 356 342
rect 358 340 359 342
rect 325 338 339 339
rect 355 338 359 340
rect 321 337 339 338
rect 328 330 332 332
rect 328 328 329 330
rect 331 328 332 330
rect 328 318 332 328
rect 335 326 339 337
rect 370 342 374 346
rect 370 338 390 342
rect 386 335 390 338
rect 378 333 382 335
rect 378 331 379 333
rect 381 331 382 333
rect 378 326 382 331
rect 386 333 392 335
rect 386 331 389 333
rect 391 331 392 333
rect 386 329 392 331
rect 335 322 342 326
rect 338 321 342 322
rect 338 319 339 321
rect 341 319 342 321
rect 328 314 334 318
rect 338 317 342 319
rect 386 318 390 329
rect 350 317 390 318
rect 350 315 374 317
rect 376 315 390 317
rect 350 314 390 315
rect 330 310 354 314
rect 373 310 377 314
rect 425 349 431 356
rect 425 347 427 349
rect 429 347 431 349
rect 425 346 431 347
rect 436 347 440 349
rect 436 345 437 347
rect 439 345 440 347
rect 436 343 440 345
rect 445 347 451 356
rect 479 354 481 356
rect 483 354 485 356
rect 479 353 485 354
rect 537 353 541 356
rect 580 354 582 356
rect 584 354 586 356
rect 580 353 586 354
rect 638 353 642 356
rect 679 354 681 356
rect 683 354 685 356
rect 679 353 685 354
rect 737 353 741 356
rect 537 351 538 353
rect 540 351 541 353
rect 638 351 639 353
rect 641 351 642 353
rect 737 351 738 353
rect 740 351 741 353
rect 507 350 532 351
rect 445 345 447 347
rect 449 345 451 347
rect 445 344 451 345
rect 492 349 502 350
rect 492 347 498 349
rect 500 347 502 349
rect 492 346 502 347
rect 507 349 528 350
rect 507 347 508 349
rect 510 348 528 349
rect 530 348 532 350
rect 537 349 541 351
rect 608 350 633 351
rect 510 347 532 348
rect 423 339 440 343
rect 423 333 427 339
rect 423 331 424 333
rect 426 331 427 333
rect 423 318 427 331
rect 446 319 447 335
rect 419 311 420 317
rect 423 314 435 318
rect 360 309 366 310
rect 360 307 362 309
rect 364 307 366 309
rect 246 300 248 302
rect 250 300 252 302
rect 281 302 287 303
rect 281 300 283 302
rect 285 300 287 302
rect 325 302 331 303
rect 325 300 327 302
rect 329 300 331 302
rect 360 302 366 307
rect 373 308 374 310
rect 376 308 377 310
rect 373 306 377 308
rect 382 309 388 310
rect 382 307 384 309
rect 386 307 388 309
rect 360 300 362 302
rect 364 300 366 302
rect 382 302 388 307
rect 431 309 435 314
rect 492 342 496 346
rect 476 338 496 342
rect 476 335 480 338
rect 474 333 480 335
rect 474 331 475 333
rect 477 331 480 333
rect 474 329 480 331
rect 476 318 480 329
rect 484 333 488 335
rect 507 342 511 347
rect 507 340 508 342
rect 510 340 511 342
rect 507 338 511 340
rect 516 342 531 343
rect 516 340 518 342
rect 520 341 531 342
rect 520 340 545 341
rect 516 339 541 340
rect 527 338 541 339
rect 543 338 545 340
rect 527 337 545 338
rect 484 331 485 333
rect 487 331 488 333
rect 484 326 488 331
rect 527 326 531 337
rect 524 322 531 326
rect 534 330 538 332
rect 534 328 535 330
rect 537 328 538 330
rect 524 321 528 322
rect 524 319 525 321
rect 527 319 528 321
rect 476 317 516 318
rect 524 317 528 319
rect 534 318 538 328
rect 476 315 490 317
rect 492 315 516 317
rect 476 314 516 315
rect 532 314 538 318
rect 489 310 493 314
rect 512 310 536 314
rect 593 349 603 350
rect 593 347 599 349
rect 601 347 603 349
rect 593 346 603 347
rect 608 349 629 350
rect 608 347 609 349
rect 611 348 629 349
rect 631 348 633 350
rect 638 349 642 351
rect 707 350 732 351
rect 611 347 633 348
rect 593 342 597 346
rect 577 338 597 342
rect 577 335 581 338
rect 575 333 581 335
rect 575 331 576 333
rect 578 331 581 333
rect 575 329 581 331
rect 577 318 581 329
rect 585 333 589 335
rect 608 342 612 347
rect 608 340 609 342
rect 611 340 612 342
rect 608 338 612 340
rect 617 342 632 343
rect 617 340 619 342
rect 621 341 632 342
rect 621 340 646 341
rect 617 339 642 340
rect 628 338 642 339
rect 644 338 646 340
rect 628 337 646 338
rect 585 331 586 333
rect 588 331 589 333
rect 585 326 589 331
rect 628 326 632 337
rect 625 322 632 326
rect 635 330 639 332
rect 635 328 636 330
rect 638 328 639 330
rect 625 321 629 322
rect 625 319 626 321
rect 628 319 629 321
rect 577 317 617 318
rect 625 317 629 319
rect 635 318 639 328
rect 577 315 591 317
rect 593 315 617 317
rect 577 314 617 315
rect 633 314 639 318
rect 590 310 594 314
rect 613 310 637 314
rect 692 349 702 350
rect 692 347 698 349
rect 700 347 702 349
rect 692 346 702 347
rect 707 349 728 350
rect 707 347 708 349
rect 710 348 728 349
rect 730 348 732 350
rect 737 349 741 351
rect 710 347 732 348
rect 692 342 696 346
rect 676 338 696 342
rect 676 335 680 338
rect 674 333 680 335
rect 674 331 675 333
rect 677 331 680 333
rect 674 329 680 331
rect 676 318 680 329
rect 684 333 688 335
rect 707 342 711 347
rect 707 340 708 342
rect 710 340 711 342
rect 707 338 711 340
rect 716 342 731 343
rect 716 340 718 342
rect 720 341 731 342
rect 720 340 745 341
rect 716 339 741 340
rect 727 338 741 339
rect 743 338 745 340
rect 727 337 745 338
rect 684 331 685 333
rect 687 331 688 333
rect 684 326 688 331
rect 727 326 731 337
rect 724 322 731 326
rect 734 330 738 332
rect 734 328 735 330
rect 737 328 738 330
rect 724 321 728 322
rect 724 319 725 321
rect 727 319 728 321
rect 676 317 716 318
rect 724 317 728 319
rect 734 318 738 328
rect 676 315 690 317
rect 692 315 716 317
rect 676 314 716 315
rect 732 314 738 318
rect 689 310 693 314
rect 712 310 736 314
rect 478 309 484 310
rect 431 308 451 309
rect 431 306 447 308
rect 449 306 451 308
rect 431 305 451 306
rect 478 307 480 309
rect 482 307 484 309
rect 382 300 384 302
rect 386 300 388 302
rect 478 302 484 307
rect 489 308 490 310
rect 492 308 493 310
rect 489 306 493 308
rect 500 309 506 310
rect 500 307 502 309
rect 504 307 506 309
rect 478 300 480 302
rect 482 300 484 302
rect 500 302 506 307
rect 579 309 585 310
rect 579 307 581 309
rect 583 307 585 309
rect 500 300 502 302
rect 504 300 506 302
rect 535 302 541 303
rect 535 300 537 302
rect 539 300 541 302
rect 579 302 585 307
rect 590 308 591 310
rect 593 308 594 310
rect 590 306 594 308
rect 601 309 607 310
rect 601 307 603 309
rect 605 307 607 309
rect 579 300 581 302
rect 583 300 585 302
rect 601 302 607 307
rect 678 309 684 310
rect 678 307 680 309
rect 682 307 684 309
rect 601 300 603 302
rect 605 300 607 302
rect 636 302 642 303
rect 636 300 638 302
rect 640 300 642 302
rect 678 302 684 307
rect 689 308 690 310
rect 692 308 693 310
rect 689 306 693 308
rect 700 309 706 310
rect 700 307 702 309
rect 704 307 706 309
rect 678 300 680 302
rect 682 300 684 302
rect 700 302 706 307
rect 700 300 702 302
rect 704 300 706 302
rect 735 302 741 303
rect 735 300 737 302
rect 739 300 741 302
rect 122 282 124 284
rect 126 282 128 284
rect 87 278 107 279
rect 87 276 103 278
rect 105 276 107 278
rect 87 275 107 276
rect 122 277 128 282
rect 144 282 146 284
rect 148 282 150 284
rect 122 275 124 277
rect 126 275 128 277
rect 75 267 76 273
rect 87 270 91 275
rect 122 274 128 275
rect 133 276 137 278
rect 133 274 134 276
rect 136 274 137 276
rect 144 277 150 282
rect 179 282 181 284
rect 183 282 185 284
rect 179 281 185 282
rect 223 282 225 284
rect 227 282 229 284
rect 144 275 146 277
rect 148 275 150 277
rect 144 274 150 275
rect 223 277 229 282
rect 245 282 247 284
rect 249 282 251 284
rect 223 275 225 277
rect 227 275 229 277
rect 223 274 229 275
rect 234 276 238 278
rect 234 274 235 276
rect 237 274 238 276
rect 245 277 251 282
rect 280 282 282 284
rect 284 282 286 284
rect 280 281 286 282
rect 324 282 326 284
rect 328 282 330 284
rect 245 275 247 277
rect 249 275 251 277
rect 245 274 251 275
rect 324 277 330 282
rect 346 282 348 284
rect 350 282 352 284
rect 324 275 326 277
rect 328 275 330 277
rect 324 274 330 275
rect 335 276 339 278
rect 335 274 336 276
rect 338 274 339 276
rect 346 277 352 282
rect 381 282 383 284
rect 385 282 387 284
rect 381 281 387 282
rect 477 282 479 284
rect 481 282 483 284
rect 346 275 348 277
rect 350 275 352 277
rect 346 274 352 275
rect 79 266 91 270
rect 133 270 137 274
rect 156 270 180 274
rect 79 253 83 266
rect 79 251 80 253
rect 82 251 83 253
rect 79 245 83 251
rect 102 249 103 265
rect 120 269 160 270
rect 120 267 134 269
rect 136 267 160 269
rect 120 266 160 267
rect 79 241 96 245
rect 92 239 96 241
rect 81 237 87 238
rect 81 235 83 237
rect 85 235 87 237
rect 92 237 93 239
rect 95 237 96 239
rect 92 235 96 237
rect 101 239 107 240
rect 101 237 103 239
rect 105 237 107 239
rect 81 228 87 235
rect 101 228 107 237
rect 120 255 124 266
rect 168 265 172 267
rect 176 266 182 270
rect 168 263 169 265
rect 171 263 172 265
rect 168 262 172 263
rect 168 258 175 262
rect 118 253 124 255
rect 118 251 119 253
rect 121 251 124 253
rect 118 249 124 251
rect 128 253 132 258
rect 128 251 129 253
rect 131 251 132 253
rect 128 249 132 251
rect 120 246 124 249
rect 120 242 140 246
rect 136 238 140 242
rect 171 247 175 258
rect 178 256 182 266
rect 178 254 179 256
rect 181 254 182 256
rect 178 252 182 254
rect 171 246 189 247
rect 151 244 155 246
rect 171 245 185 246
rect 151 242 152 244
rect 154 242 155 244
rect 136 237 146 238
rect 136 235 142 237
rect 144 235 146 237
rect 136 234 146 235
rect 151 237 155 242
rect 160 244 185 245
rect 187 244 189 246
rect 160 242 162 244
rect 164 243 189 244
rect 164 242 175 243
rect 160 241 175 242
rect 151 235 152 237
rect 154 236 176 237
rect 154 235 172 236
rect 151 234 172 235
rect 174 234 176 236
rect 151 233 176 234
rect 181 233 185 235
rect 234 270 238 274
rect 257 270 281 274
rect 221 269 261 270
rect 221 267 235 269
rect 237 267 261 269
rect 221 266 261 267
rect 221 255 225 266
rect 269 265 273 267
rect 277 266 283 270
rect 269 263 270 265
rect 272 263 273 265
rect 269 262 273 263
rect 269 258 276 262
rect 219 253 225 255
rect 219 251 220 253
rect 222 251 225 253
rect 219 249 225 251
rect 229 253 233 258
rect 229 251 230 253
rect 232 251 233 253
rect 229 249 233 251
rect 221 246 225 249
rect 221 242 241 246
rect 237 238 241 242
rect 272 247 276 258
rect 279 256 283 266
rect 279 254 280 256
rect 282 254 283 256
rect 279 252 283 254
rect 272 246 290 247
rect 252 244 256 246
rect 272 245 286 246
rect 252 242 253 244
rect 255 242 256 244
rect 237 237 247 238
rect 237 235 243 237
rect 245 235 247 237
rect 237 234 247 235
rect 252 237 256 242
rect 261 244 286 245
rect 288 244 290 246
rect 261 242 263 244
rect 265 243 290 244
rect 265 242 276 243
rect 261 241 276 242
rect 252 235 253 237
rect 255 236 277 237
rect 255 235 273 236
rect 252 234 273 235
rect 275 234 277 236
rect 252 233 277 234
rect 282 233 286 235
rect 335 270 339 274
rect 358 270 382 274
rect 322 269 362 270
rect 322 267 336 269
rect 338 267 362 269
rect 322 266 362 267
rect 322 255 326 266
rect 370 265 374 267
rect 378 266 384 270
rect 370 263 371 265
rect 373 263 374 265
rect 370 262 374 263
rect 370 258 377 262
rect 320 253 326 255
rect 320 251 321 253
rect 323 251 326 253
rect 320 249 326 251
rect 330 253 334 258
rect 330 251 331 253
rect 333 251 334 253
rect 330 249 334 251
rect 322 246 326 249
rect 322 242 342 246
rect 338 238 342 242
rect 373 247 377 258
rect 380 256 384 266
rect 380 254 381 256
rect 383 254 384 256
rect 380 252 384 254
rect 373 246 391 247
rect 353 244 357 246
rect 373 245 387 246
rect 353 242 354 244
rect 356 242 357 244
rect 338 237 348 238
rect 338 235 344 237
rect 346 235 348 237
rect 338 234 348 235
rect 353 237 357 242
rect 362 244 387 245
rect 389 244 391 246
rect 362 242 364 244
rect 366 243 391 244
rect 366 242 377 243
rect 362 241 377 242
rect 353 235 354 237
rect 356 236 378 237
rect 356 235 374 236
rect 353 234 374 235
rect 376 234 378 236
rect 353 233 378 234
rect 383 233 387 235
rect 430 278 450 279
rect 430 276 446 278
rect 448 276 450 278
rect 430 275 450 276
rect 477 277 483 282
rect 499 282 501 284
rect 503 282 505 284
rect 477 275 479 277
rect 481 275 483 277
rect 418 267 419 273
rect 430 270 434 275
rect 477 274 483 275
rect 488 276 492 278
rect 488 274 489 276
rect 491 274 492 276
rect 499 277 505 282
rect 534 282 536 284
rect 538 282 540 284
rect 534 281 540 282
rect 578 282 580 284
rect 582 282 584 284
rect 499 275 501 277
rect 503 275 505 277
rect 499 274 505 275
rect 578 277 584 282
rect 600 282 602 284
rect 604 282 606 284
rect 578 275 580 277
rect 582 275 584 277
rect 578 274 584 275
rect 589 276 593 278
rect 589 274 590 276
rect 592 274 593 276
rect 600 277 606 282
rect 635 282 637 284
rect 639 282 641 284
rect 635 281 641 282
rect 677 282 679 284
rect 681 282 683 284
rect 600 275 602 277
rect 604 275 606 277
rect 600 274 606 275
rect 677 277 683 282
rect 699 282 701 284
rect 703 282 705 284
rect 677 275 679 277
rect 681 275 683 277
rect 677 274 683 275
rect 688 276 692 278
rect 688 274 689 276
rect 691 274 692 276
rect 699 277 705 282
rect 734 282 736 284
rect 738 282 740 284
rect 734 281 740 282
rect 699 275 701 277
rect 703 275 705 277
rect 699 274 705 275
rect 422 266 434 270
rect 488 270 492 274
rect 511 270 535 274
rect 422 253 426 266
rect 422 251 423 253
rect 425 251 426 253
rect 422 245 426 251
rect 445 249 446 265
rect 475 269 515 270
rect 475 267 489 269
rect 491 267 515 269
rect 475 266 515 267
rect 422 241 439 245
rect 435 239 439 241
rect 424 237 430 238
rect 424 235 426 237
rect 428 235 430 237
rect 435 237 436 239
rect 438 237 439 239
rect 435 235 439 237
rect 444 239 450 240
rect 444 237 446 239
rect 448 237 450 239
rect 181 231 182 233
rect 184 231 185 233
rect 282 231 283 233
rect 285 231 286 233
rect 383 231 384 233
rect 386 231 387 233
rect 123 230 129 231
rect 123 228 125 230
rect 127 228 129 230
rect 181 228 185 231
rect 224 230 230 231
rect 224 228 226 230
rect 228 228 230 230
rect 282 228 286 231
rect 325 230 331 231
rect 325 228 327 230
rect 329 228 331 230
rect 383 228 387 231
rect 424 228 430 235
rect 444 228 450 237
rect 475 255 479 266
rect 523 265 527 267
rect 531 266 537 270
rect 523 263 524 265
rect 526 263 527 265
rect 523 262 527 263
rect 523 258 530 262
rect 473 253 479 255
rect 473 251 474 253
rect 476 251 479 253
rect 473 249 479 251
rect 483 253 487 258
rect 483 251 484 253
rect 486 251 487 253
rect 483 249 487 251
rect 475 246 479 249
rect 475 242 495 246
rect 491 238 495 242
rect 526 247 530 258
rect 533 256 537 266
rect 533 254 534 256
rect 536 254 537 256
rect 533 252 537 254
rect 526 246 544 247
rect 506 244 510 246
rect 526 245 540 246
rect 506 242 507 244
rect 509 242 510 244
rect 491 237 501 238
rect 491 235 497 237
rect 499 235 501 237
rect 491 234 501 235
rect 506 237 510 242
rect 515 244 540 245
rect 542 244 544 246
rect 515 242 517 244
rect 519 243 544 244
rect 519 242 530 243
rect 515 241 530 242
rect 506 235 507 237
rect 509 236 531 237
rect 509 235 527 236
rect 506 234 527 235
rect 529 234 531 236
rect 506 233 531 234
rect 536 233 540 235
rect 589 270 593 274
rect 612 270 636 274
rect 576 269 616 270
rect 576 267 590 269
rect 592 267 616 269
rect 576 266 616 267
rect 576 255 580 266
rect 624 265 628 267
rect 632 266 638 270
rect 624 263 625 265
rect 627 263 628 265
rect 624 262 628 263
rect 624 258 631 262
rect 574 253 580 255
rect 574 251 575 253
rect 577 251 580 253
rect 574 249 580 251
rect 584 253 588 258
rect 584 251 585 253
rect 587 251 588 253
rect 584 249 588 251
rect 576 246 580 249
rect 576 242 596 246
rect 592 238 596 242
rect 627 247 631 258
rect 634 256 638 266
rect 634 254 635 256
rect 637 254 638 256
rect 634 252 638 254
rect 627 246 645 247
rect 607 244 611 246
rect 627 245 641 246
rect 607 242 608 244
rect 610 242 611 244
rect 592 237 602 238
rect 592 235 598 237
rect 600 235 602 237
rect 592 234 602 235
rect 607 237 611 242
rect 616 244 641 245
rect 643 244 645 246
rect 616 242 618 244
rect 620 243 645 244
rect 620 242 631 243
rect 616 241 631 242
rect 607 235 608 237
rect 610 236 632 237
rect 610 235 628 236
rect 607 234 628 235
rect 630 234 632 236
rect 607 233 632 234
rect 637 233 641 235
rect 688 270 692 274
rect 711 270 735 274
rect 675 269 715 270
rect 675 267 689 269
rect 691 267 715 269
rect 675 266 715 267
rect 675 255 679 266
rect 723 265 727 267
rect 731 266 737 270
rect 723 263 724 265
rect 726 263 727 265
rect 723 262 727 263
rect 723 258 730 262
rect 673 253 679 255
rect 673 251 674 253
rect 676 251 679 253
rect 673 249 679 251
rect 683 253 687 258
rect 683 251 684 253
rect 686 251 687 253
rect 683 249 687 251
rect 675 246 679 249
rect 675 242 695 246
rect 691 238 695 242
rect 726 247 730 258
rect 733 256 737 266
rect 733 254 734 256
rect 736 254 737 256
rect 733 252 737 254
rect 726 246 744 247
rect 706 244 710 246
rect 726 245 740 246
rect 706 242 707 244
rect 709 242 710 244
rect 691 237 701 238
rect 691 235 697 237
rect 699 235 701 237
rect 691 234 701 235
rect 706 237 710 242
rect 715 244 740 245
rect 742 244 744 246
rect 715 242 717 244
rect 719 243 744 244
rect 719 242 730 243
rect 715 241 730 242
rect 706 235 707 237
rect 709 236 731 237
rect 709 235 727 236
rect 706 234 727 235
rect 729 234 731 236
rect 706 233 731 234
rect 736 233 740 235
rect 536 231 537 233
rect 539 231 540 233
rect 637 231 638 233
rect 640 231 641 233
rect 736 231 737 233
rect 739 231 740 233
rect 478 230 484 231
rect 478 228 480 230
rect 482 228 484 230
rect 536 228 540 231
rect 579 230 585 231
rect 579 228 581 230
rect 583 228 585 230
rect 637 228 641 231
rect 678 230 684 231
rect 678 228 680 230
rect 682 228 684 230
rect 736 228 740 231
<< via1 >>
rect 403 579 405 581
rect 449 579 451 581
rect 494 579 496 581
rect 567 579 569 581
rect 68 575 70 577
rect 108 576 110 578
rect 146 575 148 577
rect 217 575 219 577
rect 282 575 284 577
rect 335 575 337 577
rect 370 575 372 577
rect 632 575 634 577
rect 753 576 755 578
rect 103 563 105 565
rect 81 547 83 549
rect 79 530 81 532
rect 112 547 114 549
rect 119 530 121 532
rect 143 522 145 524
rect 168 547 170 549
rect 185 530 187 532
rect 170 523 172 525
rect 232 523 234 525
rect 314 547 316 549
rect 297 530 299 532
rect 250 523 252 525
rect 312 523 314 525
rect 379 563 381 565
rect 370 547 372 549
rect 339 522 341 524
rect 363 530 365 532
rect 401 547 403 549
rect 403 530 405 532
rect 484 547 486 549
rect 467 530 469 532
rect 420 523 422 525
rect 482 523 484 525
rect 549 563 551 565
rect 540 547 542 549
rect 619 563 621 565
rect 509 522 511 524
rect 533 530 535 532
rect 571 547 573 549
rect 597 547 599 549
rect 573 530 575 532
rect 595 530 597 532
rect 628 547 630 549
rect 635 530 637 532
rect 659 522 661 524
rect 684 547 686 549
rect 701 530 703 532
rect 686 523 688 525
rect 68 507 70 509
rect 129 507 131 509
rect 193 507 195 509
rect 257 507 259 509
rect 320 507 322 509
rect 355 507 357 509
rect 387 507 389 509
rect 428 507 430 509
rect 459 507 461 509
rect 516 507 518 509
rect 606 507 608 509
rect 709 507 711 509
rect 753 507 755 509
rect 79 484 81 486
rect 81 467 83 469
rect 104 475 106 477
rect 119 484 121 486
rect 143 492 145 494
rect 112 467 114 469
rect 154 459 156 461
rect 176 475 178 477
rect 168 467 170 469
rect 232 456 234 458
rect 306 475 308 477
rect 314 467 316 469
rect 328 459 330 461
rect 250 456 252 458
rect 339 492 341 494
rect 363 484 365 486
rect 370 467 372 469
rect 403 484 405 486
rect 401 467 403 469
rect 379 454 381 456
rect 420 463 422 465
rect 500 483 502 485
rect 476 475 478 477
rect 484 467 486 469
rect 509 492 511 494
rect 533 484 535 486
rect 573 484 575 486
rect 548 475 550 477
rect 540 467 542 469
rect 595 484 597 486
rect 571 467 573 469
rect 597 467 599 469
rect 635 484 637 486
rect 659 492 661 494
rect 628 467 630 469
rect 670 459 672 461
rect 692 475 694 477
rect 684 467 686 469
rect 740 451 742 453
rect 68 434 70 436
rect 108 435 110 437
rect 146 435 148 437
rect 217 435 219 437
rect 282 435 284 437
rect 335 435 337 437
rect 370 434 372 436
rect 402 434 404 436
rect 449 435 451 437
rect 494 435 496 437
rect 753 436 755 438
rect 567 434 569 436
rect 632 434 634 436
rect 193 419 195 421
rect 93 394 95 396
rect 73 379 75 381
rect 162 403 164 405
rect 145 386 147 388
rect 250 403 252 405
rect 247 395 249 397
rect 215 379 217 381
rect 293 379 295 381
rect 331 403 333 405
rect 348 386 350 388
rect 395 379 397 381
rect 416 395 418 397
rect 439 394 441 396
rect 484 403 486 405
rect 502 395 504 397
rect 545 378 547 380
rect 585 403 587 405
rect 569 386 571 388
rect 650 394 652 396
rect 602 386 604 388
rect 684 403 686 405
rect 692 395 694 397
rect 668 386 670 388
rect 748 379 750 381
rect 65 363 67 365
rect 129 362 131 364
rect 193 363 195 365
rect 257 363 259 365
rect 320 363 322 365
rect 356 363 358 365
rect 387 363 389 365
rect 428 362 430 364
rect 459 362 461 364
rect 516 362 518 364
rect 606 363 608 365
rect 709 363 711 365
rect 753 363 755 365
rect 91 347 93 349
rect 153 347 155 349
rect 106 339 108 341
rect 123 323 125 325
rect 163 340 165 342
rect 247 340 249 342
rect 185 332 187 334
rect 295 339 297 341
rect 267 331 269 333
rect 378 347 380 349
rect 363 339 365 341
rect 380 323 382 325
rect 416 323 418 325
rect 439 332 441 334
rect 324 307 326 309
rect 502 331 504 333
rect 518 323 520 325
rect 569 340 571 342
rect 602 340 604 342
rect 650 332 652 334
rect 619 324 621 326
rect 668 340 670 342
rect 701 340 703 342
rect 718 323 720 325
rect 65 291 67 293
rect 109 292 111 294
rect 146 291 148 293
rect 217 291 219 293
rect 282 291 284 293
rect 335 291 337 293
rect 370 290 372 292
rect 403 291 405 293
rect 449 291 451 293
rect 494 291 496 293
rect 567 290 569 292
rect 632 290 634 292
rect 752 291 754 293
rect 95 250 97 252
rect 128 259 130 261
rect 146 251 148 253
rect 229 259 231 261
rect 213 242 215 244
rect 294 250 296 252
rect 246 242 248 244
rect 330 259 332 261
rect 314 242 316 244
rect 347 247 349 249
rect 415 247 417 249
rect 438 250 440 252
rect 483 259 485 261
rect 501 251 503 253
rect 584 259 586 261
rect 568 242 570 244
rect 649 250 651 252
rect 601 242 603 244
rect 683 259 685 261
rect 691 251 693 253
rect 667 242 669 244
rect 68 223 70 225
rect 709 223 711 225
rect 752 223 754 225
rect 129 218 131 220
rect 193 218 195 220
rect 257 218 259 220
rect 320 218 322 220
rect 356 218 358 220
rect 387 218 389 220
rect 428 218 430 220
rect 459 218 461 220
rect 516 218 518 220
rect 606 218 608 220
<< via2 >>
rect 403 579 405 581
rect 449 579 451 581
rect 494 579 496 581
rect 567 579 569 581
rect 68 575 70 577
rect 108 576 110 578
rect 146 575 148 577
rect 217 575 219 577
rect 282 575 284 577
rect 335 575 337 577
rect 370 575 372 577
rect 632 575 634 577
rect 753 576 755 578
rect 401 571 403 573
rect 597 571 599 573
rect 168 563 170 565
rect 314 563 316 565
rect 484 563 486 565
rect 684 563 686 565
rect 112 555 114 557
rect 540 555 542 557
rect 112 547 114 549
rect 168 547 170 549
rect 314 547 316 549
rect 401 547 403 549
rect 484 547 486 549
rect 540 547 542 549
rect 597 547 599 549
rect 684 547 686 549
rect 79 539 81 541
rect 403 539 405 541
rect 533 538 535 540
rect 635 538 637 540
rect 79 530 81 532
rect 119 530 121 532
rect 185 530 187 532
rect 297 530 299 532
rect 363 530 365 532
rect 403 530 405 532
rect 467 530 469 532
rect 533 530 535 532
rect 573 530 575 532
rect 595 530 597 532
rect 635 530 637 532
rect 701 530 703 532
rect 147 522 149 524
rect 170 523 172 525
rect 237 523 239 525
rect 250 523 252 525
rect 312 523 314 525
rect 335 522 337 524
rect 420 523 422 525
rect 482 523 484 525
rect 505 522 507 524
rect 663 522 665 524
rect 686 523 688 525
rect 68 507 70 509
rect 129 507 131 509
rect 193 507 195 509
rect 257 507 259 509
rect 320 507 322 509
rect 355 507 357 509
rect 387 507 389 509
rect 428 507 430 509
rect 459 507 461 509
rect 516 507 518 509
rect 606 507 608 509
rect 709 507 711 509
rect 753 507 755 509
rect 185 492 187 494
rect 297 492 299 494
rect 467 492 469 494
rect 701 492 703 494
rect 79 484 81 486
rect 119 484 121 486
rect 363 484 365 486
rect 403 484 405 486
rect 459 483 461 485
rect 533 484 535 486
rect 573 484 575 486
rect 595 484 597 486
rect 635 484 637 486
rect 100 475 102 477
rect 170 475 172 477
rect 249 475 251 477
rect 298 475 300 477
rect 312 475 314 477
rect 482 475 484 477
rect 559 475 561 477
rect 686 475 688 477
rect 108 467 110 469
rect 147 467 149 469
rect 209 467 211 469
rect 259 467 261 469
rect 335 467 337 469
rect 401 467 403 469
rect 505 467 507 469
rect 540 467 542 469
rect 597 467 599 469
rect 663 467 665 469
rect 410 463 412 465
rect 154 459 156 461
rect 259 459 261 461
rect 228 456 230 458
rect 654 459 656 461
rect 250 456 252 458
rect 379 454 381 456
rect 401 454 403 456
rect 597 454 599 456
rect 740 451 742 453
rect 108 446 110 448
rect 540 446 542 448
rect 68 434 70 436
rect 108 435 110 437
rect 146 435 148 437
rect 217 435 219 437
rect 282 435 284 437
rect 335 435 337 437
rect 370 434 372 436
rect 402 434 404 436
rect 449 435 451 437
rect 494 435 496 437
rect 567 434 569 436
rect 632 434 634 436
rect 753 436 755 438
rect 331 419 333 421
rect 379 419 381 421
rect 684 419 686 421
rect 298 411 300 413
rect 484 411 486 413
rect 559 411 561 413
rect 692 411 694 413
rect 201 403 203 405
rect 250 403 252 405
rect 331 403 333 405
rect 359 403 361 405
rect 459 403 461 405
rect 484 403 486 405
rect 585 403 587 405
rect 684 403 686 405
rect 93 394 95 396
rect 154 394 156 396
rect 162 394 164 396
rect 692 395 694 397
rect 153 386 155 388
rect 201 387 203 389
rect 305 387 307 389
rect 348 386 350 388
rect 73 379 75 381
rect 185 379 187 381
rect 247 379 249 381
rect 305 378 307 380
rect 359 378 361 380
rect 395 379 397 381
rect 545 378 547 380
rect 701 379 703 381
rect 420 370 422 372
rect 585 370 587 372
rect 65 363 67 365
rect 129 362 131 364
rect 193 363 195 365
rect 257 363 259 365
rect 320 363 322 365
rect 356 363 358 365
rect 387 363 389 365
rect 428 362 430 364
rect 459 362 461 364
rect 516 362 518 364
rect 606 363 608 365
rect 709 363 711 365
rect 753 363 755 365
rect 91 347 93 349
rect 153 347 155 349
rect 348 347 350 349
rect 247 340 249 342
rect 701 340 703 342
rect 185 332 187 334
rect 410 331 412 333
rect 209 323 211 325
rect 545 323 547 325
rect 654 324 656 326
rect 740 323 742 325
rect 324 307 326 309
rect 324 299 326 301
rect 691 299 693 301
rect 65 291 67 293
rect 109 292 111 294
rect 146 291 148 293
rect 217 291 219 293
rect 282 291 284 293
rect 335 291 337 293
rect 370 290 372 292
rect 403 291 405 293
rect 449 291 451 293
rect 494 291 496 293
rect 567 290 569 292
rect 632 290 634 292
rect 752 291 754 293
rect 395 281 397 283
rect 483 281 485 283
rect 228 267 230 269
rect 330 267 332 269
rect 73 259 75 261
rect 162 259 164 261
rect 330 259 332 261
rect 483 259 485 261
rect 584 259 586 261
rect 683 259 685 261
rect 691 251 693 253
rect 237 234 239 236
rect 584 234 586 236
rect 101 226 103 228
rect 683 226 685 228
rect 68 223 70 225
rect 709 223 711 225
rect 752 223 754 225
rect 129 218 131 220
rect 193 218 195 220
rect 257 218 259 220
rect 320 218 322 220
rect 356 218 358 220
rect 387 218 389 220
rect 428 218 430 220
rect 459 218 461 220
rect 516 218 518 220
rect 606 218 608 220
<< via3 >>
rect 403 579 405 581
rect 449 579 451 581
rect 494 579 496 581
rect 567 579 569 581
rect 68 575 70 577
rect 108 576 110 578
rect 146 575 148 577
rect 217 575 219 577
rect 282 575 284 577
rect 335 575 337 577
rect 370 575 372 577
rect 632 575 634 577
rect 753 576 755 578
rect 68 507 70 509
rect 129 507 131 509
rect 68 434 70 436
rect 193 507 195 509
rect 108 435 110 437
rect 146 435 148 437
rect 65 363 67 365
rect 65 291 67 293
rect 129 362 131 364
rect 109 292 111 294
rect 146 291 148 293
rect 193 363 195 365
rect 217 435 219 437
rect 217 291 219 293
rect 257 507 259 509
rect 282 435 284 437
rect 320 507 322 509
rect 355 507 357 509
rect 387 507 389 509
rect 335 435 337 437
rect 370 434 372 436
rect 402 434 404 436
rect 257 363 259 365
rect 320 363 322 365
rect 356 363 358 365
rect 387 363 389 365
rect 282 291 284 293
rect 335 291 337 293
rect 370 290 372 292
rect 428 507 430 509
rect 459 507 461 509
rect 449 435 451 437
rect 516 507 518 509
rect 606 507 608 509
rect 494 435 496 437
rect 709 507 711 509
rect 753 507 755 509
rect 567 434 569 436
rect 632 434 634 436
rect 428 362 430 364
rect 459 362 461 364
rect 516 362 518 364
rect 606 363 608 365
rect 709 363 711 365
rect 753 436 755 438
rect 753 363 755 365
rect 403 291 405 293
rect 449 291 451 293
rect 494 291 496 293
rect 567 290 569 292
rect 632 290 634 292
rect 752 291 754 293
rect 68 223 70 225
rect 709 223 711 225
rect 752 223 754 225
rect 129 218 131 220
rect 193 218 195 220
rect 257 218 259 220
rect 320 218 322 220
rect 356 218 358 220
rect 387 218 389 220
rect 428 218 430 220
rect 459 218 461 220
rect 516 218 518 220
rect 606 218 608 220
<< via4 >>
rect 129 598 131 600
rect 49 507 51 509
rect 49 363 51 365
rect 49 223 51 225
rect 108 590 110 592
rect 57 575 59 577
rect 68 575 70 577
rect 68 507 70 509
rect 57 434 59 436
rect 68 434 70 436
rect 65 363 67 365
rect 193 598 195 600
rect 57 291 59 293
rect 65 291 67 293
rect 68 223 70 225
rect 108 208 110 210
rect 146 590 148 592
rect 146 208 148 210
rect 257 598 259 600
rect 129 200 131 202
rect 217 590 219 592
rect 217 208 219 210
rect 320 598 322 600
rect 193 200 195 202
rect 282 590 284 592
rect 282 208 284 210
rect 356 598 358 600
rect 257 200 259 202
rect 335 590 337 592
rect 387 598 389 600
rect 335 208 337 210
rect 320 200 322 202
rect 370 590 372 592
rect 370 208 372 210
rect 428 598 430 600
rect 403 590 405 592
rect 356 200 358 202
rect 403 208 405 210
rect 459 598 461 600
rect 387 200 389 202
rect 449 590 451 592
rect 449 208 451 210
rect 516 598 518 600
rect 428 200 430 202
rect 494 590 496 592
rect 494 208 496 210
rect 606 598 608 600
rect 459 200 461 202
rect 567 590 569 592
rect 567 208 569 210
rect 709 598 711 600
rect 516 200 518 202
rect 632 590 634 592
rect 632 208 634 210
rect 753 576 755 578
rect 763 576 765 578
rect 753 507 755 509
rect 753 436 755 438
rect 763 436 765 438
rect 753 363 755 365
rect 752 291 754 293
rect 763 291 765 293
rect 606 200 608 202
rect 752 223 754 225
rect 771 507 773 509
rect 771 363 773 365
rect 771 223 773 225
rect 709 200 711 202
<< labels >>
rlabel alu1 153 475 153 475 1 p3
rlabel alu1 154 464 154 464 1 p3
rlabel alu1 226 452 226 452 1 p2
rlabel alu1 234 476 234 476 1 p2
rlabel alu1 226 564 226 564 1 p1
rlabel alu1 234 540 234 540 1 p1
rlabel alu1 190 576 190 576 4 vdd
rlabel alu1 190 512 190 512 4 vss
rlabel alu1 190 504 190 504 2 vss
rlabel alu1 121 468 121 468 1 b2
rlabel alu1 113 460 113 460 1 b2
rlabel alu1 129 540 129 540 1 a3
rlabel alu1 121 536 121 536 1 a3
rlabel alu1 121 548 121 548 1 b3
rlabel alu1 113 556 113 556 1 b3
rlabel alu1 129 504 129 504 2 vss
rlabel alu1 129 576 129 576 4 vdd
rlabel alu1 129 512 129 512 4 vss
rlabel alu1 105 472 105 472 1 p0
rlabel alu1 97 492 97 492 1 p0
rlabel alu1 73 556 73 556 1 b3
rlabel alu1 81 548 81 548 1 b3
rlabel alu1 89 540 89 540 1 a2
rlabel alu1 81 536 81 536 1 a2
rlabel alu1 73 460 73 460 1 b2
rlabel alu1 81 468 81 468 1 b2
rlabel alu1 89 476 89 476 1 a2
rlabel alu1 81 480 81 480 1 a2
rlabel alu1 89 504 89 504 2 vss
rlabel alu1 89 576 89 576 4 vdd
rlabel alu1 89 512 89 512 4 vss
rlabel alu1 120 480 120 480 1 a3
rlabel alu1 363 480 363 480 1 a3
rlabel alu1 363 536 363 536 1 a3
rlabel alu1 363 548 363 548 1 b1
rlabel alu1 371 556 371 556 1 b1
rlabel alu1 411 556 411 556 1 b1
rlabel via1 403 548 403 548 1 b1
rlabel alu1 371 460 371 460 1 b0
rlabel alu1 363 468 363 468 1 b0
rlabel via1 403 468 403 468 1 b0
rlabel alu1 411 460 411 460 1 b0
rlabel alu1 258 564 258 564 1 q1
rlabel alu1 250 540 250 540 1 q1
rlabel alu1 258 452 258 452 1 q2
rlabel alu1 250 476 250 476 1 q2
rlabel alu1 330 464 330 464 1 q3
rlabel alu1 331 475 331 475 1 q3
rlabel alu1 379 472 379 472 1 q0
rlabel alu1 387 492 387 492 1 q0
rlabel alu1 294 576 294 576 6 vdd
rlabel alu1 294 512 294 512 6 vss
rlabel alu1 294 504 294 504 8 vss
rlabel alu1 355 540 355 540 1 a3
rlabel alu1 355 504 355 504 8 vss
rlabel alu1 355 576 355 576 6 vdd
rlabel alu1 355 512 355 512 6 vss
rlabel alu1 395 540 395 540 1 a2
rlabel alu1 403 536 403 536 1 a2
rlabel alu1 395 476 395 476 1 a2
rlabel alu1 403 480 403 480 1 a2
rlabel alu1 395 504 395 504 8 vss
rlabel alu1 395 576 395 576 6 vdd
rlabel alu1 395 512 395 512 6 vss
rlabel alu1 533 480 533 480 1 a1
rlabel alu1 525 540 525 540 1 a1
rlabel alu1 533 536 533 536 1 a1
rlabel alu1 565 540 565 540 1 a0
rlabel alu1 573 536 573 536 1 a0
rlabel alu1 573 480 573 480 1 a0
rlabel alu1 565 476 565 476 1 a0
rlabel alu1 428 564 428 564 1 r1
rlabel alu1 420 540 420 540 1 r1
rlabel alu1 420 476 420 476 1 r2
rlabel alu1 428 452 428 452 1 r2
rlabel alu1 501 475 501 475 1 r3
rlabel alu1 500 464 500 464 1 r3
rlabel alu1 557 492 557 492 1 r0
rlabel alu1 549 472 549 472 1 r0
rlabel alu1 464 576 464 576 6 vdd
rlabel alu1 464 512 464 512 6 vss
rlabel alu1 464 504 464 504 8 vss
rlabel alu1 533 468 533 468 1 b2
rlabel alu1 541 460 541 460 1 b2
rlabel alu1 533 548 533 548 1 b3
rlabel alu1 541 556 541 556 1 b3
rlabel alu1 525 504 525 504 8 vss
rlabel alu1 525 576 525 576 6 vdd
rlabel alu1 525 512 525 512 6 vss
rlabel alu1 581 556 581 556 1 b3
rlabel alu1 573 548 573 548 1 b3
rlabel alu1 581 460 581 460 1 b2
rlabel alu1 573 468 573 468 1 b2
rlabel alu1 565 504 565 504 8 vss
rlabel alu1 565 576 565 576 6 vdd
rlabel alu1 565 512 565 512 6 vss
rlabel alu1 636 480 636 480 1 a1
rlabel alu1 645 540 645 540 1 a1
rlabel alu1 637 536 637 536 1 a1
rlabel alu1 637 548 637 548 1 b1
rlabel alu1 629 556 629 556 1 b1
rlabel alu1 589 556 589 556 1 b1
rlabel via1 597 548 597 548 1 b1
rlabel alu1 605 540 605 540 1 a0
rlabel alu1 597 536 597 536 1 a0
rlabel alu1 637 468 637 468 1 b0
rlabel alu1 629 460 629 460 1 b0
rlabel via1 597 468 597 468 1 b0
rlabel alu1 589 460 589 460 1 b0
rlabel alu1 597 480 597 480 1 a0
rlabel alu1 605 476 605 476 1 a0
rlabel alu1 742 564 742 564 1 o1
rlabel alu1 750 540 750 540 1 o1
rlabel alu1 742 452 742 452 1 s2
rlabel alu1 669 475 669 475 1 s3
rlabel alu1 670 464 670 464 1 s3
rlabel alu1 613 492 613 492 1 o0
rlabel alu1 621 472 621 472 1 o0
rlabel alu1 706 576 706 576 4 vdd
rlabel alu1 706 512 706 512 4 vss
rlabel alu1 706 504 706 504 2 vss
rlabel alu1 645 504 645 504 2 vss
rlabel alu1 645 576 645 576 4 vdd
rlabel alu1 645 512 645 512 4 vss
rlabel alu1 605 504 605 504 2 vss
rlabel alu1 605 576 605 576 4 vdd
rlabel alu1 605 512 605 512 4 vss
rlabel alu1 750 476 750 476 1 s2
rlabel alu1 749 255 749 255 1 o4
rlabel alu1 701 260 701 260 1 p0
rlabel alu1 701 248 701 248 1 u0
rlabel alu1 705 288 705 288 4 vdd
rlabel alu1 705 224 705 224 4 vss
rlabel alu1 706 368 706 368 4 vss
rlabel alu1 706 432 706 432 4 vdd
rlabel alu1 702 392 702 392 1 r0
rlabel alu1 694 396 694 396 1 r0
rlabel pmos 686 404 686 404 1 q0
rlabel alu1 694 404 694 404 1 q0
rlabel alu1 702 404 702 404 1 q0
rlabel alu1 710 404 710 404 1 q0
rlabel alu1 718 400 718 400 1 q0
rlabel alu1 706 360 706 360 2 vss
rlabel alu1 706 296 706 296 2 vdd
rlabel alu1 701 324 701 324 1 s2
rlabel alu1 711 324 711 324 1 s2
rlabel alu1 750 399 750 399 1 t5
rlabel alu1 669 333 669 333 1 t4
rlabel alu1 669 399 669 399 1 t3
rlabel alu1 681 380 681 380 1 t3
rlabel alu1 750 333 750 333 1 o2
rlabel alu1 605 324 605 324 1 s3
rlabel alu1 607 360 607 360 2 vss
rlabel alu1 607 296 607 296 2 vdd
rlabel pmos 587 404 587 404 1 r1
rlabel alu1 595 404 595 404 1 r1
rlabel alu1 603 404 603 404 1 r1
rlabel alu1 611 404 611 404 1 r1
rlabel alu1 619 400 619 400 1 r1
rlabel alu1 607 368 607 368 4 vss
rlabel alu1 607 432 607 432 4 vdd
rlabel alu1 606 288 606 288 4 vdd
rlabel alu1 606 224 606 224 4 vss
rlabel alu1 601 260 601 260 1 p1
rlabel alu1 550 325 550 325 1 o3
rlabel alu1 550 399 550 399 1 t6
rlabel alu1 506 360 506 360 2 vss
rlabel alu1 506 296 506 296 2 vdd
rlabel alu1 518 400 518 400 1 q1
rlabel alu1 510 404 510 404 1 q1
rlabel alu1 502 404 502 404 1 q1
rlabel alu1 494 404 494 404 1 q1
rlabel pmos 486 404 486 404 1 q1
rlabel alu1 506 368 506 368 4 vss
rlabel alu1 506 432 506 432 4 vdd
rlabel alu1 505 288 505 288 4 vdd
rlabel alu1 505 224 505 224 4 vss
rlabel alu1 502 260 502 260 1 u1
rlabel alu1 549 257 549 257 1 o5
rlabel alu1 417 327 417 327 1 t2
rlabel alu1 417 399 417 399 1 t1
rlabel alu1 433 296 433 296 8 vdd
rlabel alu1 433 360 433 360 8 vss
rlabel alu1 433 432 433 432 6 vdd
rlabel alu1 433 368 433 368 6 vss
rlabel alu1 432 224 432 224 6 vss
rlabel alu1 432 288 432 288 6 vdd
rlabel alu1 397 390 397 390 1 u1
rlabel alu1 316 325 316 325 1 u0
rlabel alu1 353 432 353 432 4 vdd
rlabel alu1 353 368 353 368 4 vss
rlabel alu1 360 296 360 296 8 vdd
rlabel alu1 360 360 360 360 8 vss
rlabel alu1 396 256 396 256 1 o6
rlabel alu1 348 260 348 260 1 p2
rlabel alu1 352 288 352 288 4 vdd
rlabel alu1 352 224 352 224 4 vss
rlabel alu1 256 324 256 324 1 r2
rlabel alu1 248 324 248 324 1 r2
rlabel alu1 240 324 240 324 1 r2
rlabel pmos 232 324 232 324 1 r2
rlabel alu1 263 400 263 400 1 q2
rlabel alu1 255 404 255 404 1 q2
rlabel alu1 247 404 247 404 1 q2
rlabel alu1 239 404 239 404 1 q2
rlabel pmos 231 404 231 404 1 q2
rlabel alu1 251 368 251 368 4 vss
rlabel alu1 251 432 251 432 4 vdd
rlabel alu1 252 296 252 296 2 vdd
rlabel alu1 252 360 252 360 2 vss
rlabel alu1 248 260 248 260 1 p3
rlabel alu1 251 224 251 224 4 vss
rlabel alu1 251 288 251 288 4 vdd
rlabel alu1 73 400 73 400 1 ca1
rlabel alu1 162 400 162 400 1 r3
rlabel alu1 154 404 154 404 1 r3
rlabel alu1 146 404 146 404 1 r3
rlabel alu1 138 404 138 404 1 r3
rlabel pmos 130 404 130 404 1 r3
rlabel alu1 115 324 115 324 1 q3
rlabel alu1 107 324 107 324 1 q3
rlabel alu1 99 324 99 324 1 q3
rlabel pmos 91 324 91 324 1 q3
rlabel alu1 179 296 179 296 8 vdd
rlabel alu1 179 360 179 360 8 vss
rlabel alu1 171 308 171 308 8 z
rlabel alu1 163 328 163 328 8 z
rlabel alu1 111 296 111 296 2 vdd
rlabel alu1 111 360 111 360 2 vss
rlabel alu0 122 400 122 400 4 con
rlabel alu1 150 368 150 368 4 vss
rlabel alu1 150 432 150 432 4 vdd
rlabel alu1 89 432 89 432 6 vdd
rlabel alu1 89 368 89 368 6 vss
rlabel alu1 194 256 194 256 1 o7
rlabel alu1 148 260 148 260 1 ca1
rlabel alu1 150 224 150 224 4 vss
rlabel alu1 150 288 150 288 4 vdd
rlabel alu1 89 288 89 288 6 vdd
rlabel alu1 89 224 89 224 6 vss
rlabel alu1 668 248 668 248 1 x1
rlabel alu1 416 257 416 257 1 x2
rlabel alu1 315 253 315 253 1 x3
rlabel alu1 73 254 73 254 1 ca3
<< end >>
