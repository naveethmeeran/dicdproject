magic
tech scmos
timestamp 1510248381
<< ab >>
rect 29 245 69 389
rect 71 245 198 389
rect 206 245 333 389
rect 335 245 375 389
rect 376 245 503 389
rect 505 245 585 389
rect 587 245 714 389
rect 29 173 413 245
rect 27 169 413 173
rect 24 109 413 169
rect 27 101 413 109
rect 426 101 714 245
rect 29 29 69 101
rect 70 30 412 101
rect 70 29 88 30
rect 92 29 152 30
rect 156 29 216 30
rect 220 29 279 30
rect 283 29 315 30
rect 319 29 346 30
rect 350 29 387 30
rect 391 29 412 30
rect 425 30 713 101
rect 425 29 475 30
rect 479 29 565 30
rect 569 29 713 30
<< nwell >>
rect 24 349 718 394
rect 24 205 718 285
rect 24 61 718 141
<< pwell >>
rect 24 285 718 349
rect 24 141 718 205
rect 24 24 718 61
<< poly >>
rect 38 383 40 387
rect 48 383 50 387
rect 58 383 60 387
rect 78 383 80 387
rect 88 383 90 387
rect 98 383 100 387
rect 119 383 121 387
rect 129 383 131 387
rect 139 383 141 387
rect 38 360 40 364
rect 34 358 40 360
rect 34 356 36 358
rect 38 356 40 358
rect 34 354 40 356
rect 38 343 40 354
rect 48 352 50 364
rect 78 360 80 364
rect 74 358 80 360
rect 74 356 76 358
rect 78 356 80 358
rect 58 352 60 355
rect 74 354 80 356
rect 44 350 50 352
rect 44 348 46 350
rect 48 348 50 350
rect 44 346 50 348
rect 54 350 60 352
rect 54 348 56 350
rect 58 348 60 350
rect 54 346 60 348
rect 45 343 47 346
rect 58 343 60 346
rect 78 343 80 354
rect 88 352 90 364
rect 157 380 159 385
rect 164 380 166 385
rect 187 383 189 387
rect 215 383 217 387
rect 174 371 176 376
rect 238 380 240 385
rect 245 380 247 385
rect 263 383 265 387
rect 273 383 275 387
rect 283 383 285 387
rect 304 383 306 387
rect 314 383 316 387
rect 324 383 326 387
rect 344 383 346 387
rect 354 383 356 387
rect 364 383 366 387
rect 385 383 387 387
rect 228 371 230 376
rect 174 355 176 358
rect 98 352 100 355
rect 119 352 121 355
rect 129 352 131 355
rect 139 352 141 355
rect 157 352 159 355
rect 164 352 166 355
rect 174 353 183 355
rect 84 350 90 352
rect 84 348 86 350
rect 88 348 90 350
rect 84 346 90 348
rect 94 350 100 352
rect 94 348 96 350
rect 98 348 100 350
rect 94 346 100 348
rect 117 350 123 352
rect 117 348 119 350
rect 121 348 123 350
rect 117 346 123 348
rect 127 350 133 352
rect 127 348 129 350
rect 131 348 133 350
rect 127 346 133 348
rect 137 350 159 352
rect 137 348 139 350
rect 141 348 146 350
rect 148 348 159 350
rect 137 346 159 348
rect 163 350 169 352
rect 163 348 165 350
rect 167 348 169 350
rect 163 346 169 348
rect 85 343 87 346
rect 98 343 100 346
rect 38 325 40 330
rect 45 325 47 330
rect 58 324 60 329
rect 78 325 80 330
rect 85 325 87 330
rect 119 337 121 346
rect 130 343 132 346
rect 137 343 139 346
rect 157 343 159 346
rect 167 343 169 346
rect 177 351 179 353
rect 181 351 183 353
rect 177 349 183 351
rect 98 324 100 329
rect 177 336 179 349
rect 187 345 189 358
rect 183 343 189 345
rect 183 341 185 343
rect 187 341 189 343
rect 183 339 189 341
rect 187 336 189 339
rect 215 345 217 358
rect 228 355 230 358
rect 221 353 230 355
rect 221 351 223 353
rect 225 351 227 353
rect 238 352 240 355
rect 245 352 247 355
rect 263 352 265 355
rect 273 352 275 355
rect 283 352 285 355
rect 304 352 306 355
rect 314 352 316 364
rect 324 360 326 364
rect 324 358 330 360
rect 324 356 326 358
rect 328 356 330 358
rect 324 354 330 356
rect 221 349 227 351
rect 215 343 221 345
rect 215 341 217 343
rect 219 341 221 343
rect 215 339 221 341
rect 215 336 217 339
rect 225 336 227 349
rect 235 350 241 352
rect 235 348 237 350
rect 239 348 241 350
rect 235 346 241 348
rect 245 350 267 352
rect 245 348 256 350
rect 258 348 263 350
rect 265 348 267 350
rect 245 346 267 348
rect 271 350 277 352
rect 271 348 273 350
rect 275 348 277 350
rect 271 346 277 348
rect 281 350 287 352
rect 281 348 283 350
rect 285 348 287 350
rect 281 346 287 348
rect 304 350 310 352
rect 304 348 306 350
rect 308 348 310 350
rect 304 346 310 348
rect 314 350 320 352
rect 314 348 316 350
rect 318 348 320 350
rect 314 346 320 348
rect 235 343 237 346
rect 245 343 247 346
rect 265 343 267 346
rect 272 343 274 346
rect 157 324 159 329
rect 167 324 169 329
rect 119 319 121 323
rect 130 319 132 323
rect 137 319 139 323
rect 177 321 179 326
rect 187 319 189 323
rect 215 319 217 323
rect 225 321 227 326
rect 235 324 237 329
rect 245 324 247 329
rect 283 337 285 346
rect 304 343 306 346
rect 317 343 319 346
rect 324 343 326 354
rect 344 352 346 355
rect 354 352 356 364
rect 364 360 366 364
rect 364 358 370 360
rect 408 380 410 385
rect 415 380 417 385
rect 433 383 435 387
rect 443 383 445 387
rect 453 383 455 387
rect 474 383 476 387
rect 484 383 486 387
rect 494 383 496 387
rect 514 383 516 387
rect 524 383 526 387
rect 534 383 536 387
rect 554 383 556 387
rect 564 383 566 387
rect 574 383 576 387
rect 594 383 596 387
rect 604 383 606 387
rect 614 383 616 387
rect 635 383 637 387
rect 645 383 647 387
rect 655 383 657 387
rect 398 371 400 376
rect 364 356 366 358
rect 368 356 370 358
rect 364 354 370 356
rect 344 350 350 352
rect 344 348 346 350
rect 348 348 350 350
rect 344 346 350 348
rect 354 350 360 352
rect 354 348 356 350
rect 358 348 360 350
rect 354 346 360 348
rect 344 343 346 346
rect 357 343 359 346
rect 364 343 366 354
rect 385 345 387 358
rect 398 355 400 358
rect 391 353 400 355
rect 391 351 393 353
rect 395 351 397 353
rect 408 352 410 355
rect 415 352 417 355
rect 433 352 435 355
rect 443 352 445 355
rect 453 352 455 355
rect 474 352 476 355
rect 484 352 486 364
rect 494 360 496 364
rect 494 358 500 360
rect 494 356 496 358
rect 498 356 500 358
rect 494 354 500 356
rect 391 349 397 351
rect 385 343 391 345
rect 304 324 306 329
rect 317 325 319 330
rect 324 325 326 330
rect 385 341 387 343
rect 389 341 391 343
rect 385 339 391 341
rect 385 336 387 339
rect 395 336 397 349
rect 405 350 411 352
rect 405 348 407 350
rect 409 348 411 350
rect 405 346 411 348
rect 415 350 437 352
rect 415 348 426 350
rect 428 348 433 350
rect 435 348 437 350
rect 415 346 437 348
rect 441 350 447 352
rect 441 348 443 350
rect 445 348 447 350
rect 441 346 447 348
rect 451 350 457 352
rect 451 348 453 350
rect 455 348 457 350
rect 451 346 457 348
rect 474 350 480 352
rect 474 348 476 350
rect 478 348 480 350
rect 474 346 480 348
rect 484 350 490 352
rect 484 348 486 350
rect 488 348 490 350
rect 484 346 490 348
rect 405 343 407 346
rect 415 343 417 346
rect 435 343 437 346
rect 442 343 444 346
rect 344 324 346 329
rect 357 325 359 330
rect 364 325 366 330
rect 265 319 267 323
rect 272 319 274 323
rect 283 319 285 323
rect 385 319 387 323
rect 395 321 397 326
rect 405 324 407 329
rect 415 324 417 329
rect 453 337 455 346
rect 474 343 476 346
rect 487 343 489 346
rect 494 343 496 354
rect 514 352 516 355
rect 524 352 526 364
rect 534 360 536 364
rect 554 360 556 364
rect 534 358 540 360
rect 534 356 536 358
rect 538 356 540 358
rect 534 354 540 356
rect 550 358 556 360
rect 550 356 552 358
rect 554 356 556 358
rect 550 354 556 356
rect 514 350 520 352
rect 514 348 516 350
rect 518 348 520 350
rect 514 346 520 348
rect 524 350 530 352
rect 524 348 526 350
rect 528 348 530 350
rect 524 346 530 348
rect 514 343 516 346
rect 527 343 529 346
rect 534 343 536 354
rect 554 343 556 354
rect 564 352 566 364
rect 594 360 596 364
rect 590 358 596 360
rect 590 356 592 358
rect 594 356 596 358
rect 574 352 576 355
rect 590 354 596 356
rect 560 350 566 352
rect 560 348 562 350
rect 564 348 566 350
rect 560 346 566 348
rect 570 350 576 352
rect 570 348 572 350
rect 574 348 576 350
rect 570 346 576 348
rect 561 343 563 346
rect 574 343 576 346
rect 594 343 596 354
rect 604 352 606 364
rect 673 380 675 385
rect 680 380 682 385
rect 703 383 705 387
rect 690 371 692 376
rect 690 355 692 358
rect 614 352 616 355
rect 635 352 637 355
rect 645 352 647 355
rect 655 352 657 355
rect 673 352 675 355
rect 680 352 682 355
rect 690 353 699 355
rect 600 350 606 352
rect 600 348 602 350
rect 604 348 606 350
rect 600 346 606 348
rect 610 350 616 352
rect 610 348 612 350
rect 614 348 616 350
rect 610 346 616 348
rect 633 350 639 352
rect 633 348 635 350
rect 637 348 639 350
rect 633 346 639 348
rect 643 350 649 352
rect 643 348 645 350
rect 647 348 649 350
rect 643 346 649 348
rect 653 350 675 352
rect 653 348 655 350
rect 657 348 662 350
rect 664 348 675 350
rect 653 346 675 348
rect 679 350 685 352
rect 679 348 681 350
rect 683 348 685 350
rect 679 346 685 348
rect 601 343 603 346
rect 614 343 616 346
rect 474 324 476 329
rect 487 325 489 330
rect 494 325 496 330
rect 514 324 516 329
rect 527 325 529 330
rect 534 325 536 330
rect 554 325 556 330
rect 561 325 563 330
rect 435 319 437 323
rect 442 319 444 323
rect 453 319 455 323
rect 574 324 576 329
rect 594 325 596 330
rect 601 325 603 330
rect 635 337 637 346
rect 646 343 648 346
rect 653 343 655 346
rect 673 343 675 346
rect 683 343 685 346
rect 693 351 695 353
rect 697 351 699 353
rect 693 349 699 351
rect 614 324 616 329
rect 693 336 695 349
rect 703 345 705 358
rect 699 343 705 345
rect 699 341 701 343
rect 703 341 705 343
rect 699 339 705 341
rect 703 336 705 339
rect 673 324 675 329
rect 683 324 685 329
rect 635 319 637 323
rect 646 319 648 323
rect 653 319 655 323
rect 693 321 695 326
rect 703 319 705 323
rect 119 311 121 315
rect 130 311 132 315
rect 137 311 139 315
rect 38 304 40 309
rect 45 304 47 309
rect 58 305 60 310
rect 78 304 80 309
rect 85 304 87 309
rect 98 305 100 310
rect 38 280 40 291
rect 45 288 47 291
rect 58 288 60 291
rect 44 286 50 288
rect 44 284 46 286
rect 48 284 50 286
rect 44 282 50 284
rect 54 286 60 288
rect 54 284 56 286
rect 58 284 60 286
rect 54 282 60 284
rect 34 278 40 280
rect 34 276 36 278
rect 38 276 40 278
rect 34 274 40 276
rect 38 270 40 274
rect 48 270 50 282
rect 58 279 60 282
rect 78 280 80 291
rect 85 288 87 291
rect 98 288 100 291
rect 119 288 121 297
rect 157 305 159 310
rect 167 305 169 310
rect 177 308 179 313
rect 187 311 189 315
rect 215 311 217 315
rect 225 308 227 313
rect 265 311 267 315
rect 272 311 274 315
rect 283 311 285 315
rect 235 305 237 310
rect 245 305 247 310
rect 130 288 132 291
rect 137 288 139 291
rect 157 288 159 291
rect 167 288 169 291
rect 84 286 90 288
rect 84 284 86 286
rect 88 284 90 286
rect 84 282 90 284
rect 94 286 100 288
rect 94 284 96 286
rect 98 284 100 286
rect 94 282 100 284
rect 117 286 123 288
rect 117 284 119 286
rect 121 284 123 286
rect 117 282 123 284
rect 127 286 133 288
rect 127 284 129 286
rect 131 284 133 286
rect 127 282 133 284
rect 137 286 159 288
rect 137 284 139 286
rect 141 284 146 286
rect 148 284 159 286
rect 137 282 159 284
rect 163 286 169 288
rect 163 284 165 286
rect 167 284 169 286
rect 163 282 169 284
rect 177 285 179 298
rect 187 295 189 298
rect 183 293 189 295
rect 183 291 185 293
rect 187 291 189 293
rect 183 289 189 291
rect 177 283 183 285
rect 74 278 80 280
rect 74 276 76 278
rect 78 276 80 278
rect 74 274 80 276
rect 78 270 80 274
rect 88 270 90 282
rect 98 279 100 282
rect 119 279 121 282
rect 129 279 131 282
rect 139 279 141 282
rect 157 279 159 282
rect 164 279 166 282
rect 177 281 179 283
rect 181 281 183 283
rect 174 279 183 281
rect 174 276 176 279
rect 187 276 189 289
rect 215 295 217 298
rect 215 293 221 295
rect 215 291 217 293
rect 219 291 221 293
rect 215 289 221 291
rect 215 276 217 289
rect 225 285 227 298
rect 385 311 387 315
rect 304 305 306 310
rect 221 283 227 285
rect 221 281 223 283
rect 225 281 227 283
rect 235 288 237 291
rect 245 288 247 291
rect 265 288 267 291
rect 272 288 274 291
rect 283 288 285 297
rect 317 304 319 309
rect 324 304 326 309
rect 344 305 346 310
rect 357 304 359 309
rect 364 304 366 309
rect 395 308 397 313
rect 435 311 437 315
rect 442 311 444 315
rect 453 311 455 315
rect 405 305 407 310
rect 415 305 417 310
rect 385 295 387 298
rect 385 293 391 295
rect 385 291 387 293
rect 389 291 391 293
rect 304 288 306 291
rect 317 288 319 291
rect 235 286 241 288
rect 235 284 237 286
rect 239 284 241 286
rect 235 282 241 284
rect 245 286 267 288
rect 245 284 256 286
rect 258 284 263 286
rect 265 284 267 286
rect 245 282 267 284
rect 271 286 277 288
rect 271 284 273 286
rect 275 284 277 286
rect 271 282 277 284
rect 281 286 287 288
rect 281 284 283 286
rect 285 284 287 286
rect 281 282 287 284
rect 304 286 310 288
rect 304 284 306 286
rect 308 284 310 286
rect 304 282 310 284
rect 314 286 320 288
rect 314 284 316 286
rect 318 284 320 286
rect 314 282 320 284
rect 221 279 230 281
rect 238 279 240 282
rect 245 279 247 282
rect 263 279 265 282
rect 273 279 275 282
rect 283 279 285 282
rect 304 279 306 282
rect 228 276 230 279
rect 174 258 176 263
rect 38 247 40 251
rect 48 247 50 251
rect 58 247 60 251
rect 78 247 80 251
rect 88 247 90 251
rect 98 247 100 251
rect 119 247 121 251
rect 129 247 131 251
rect 139 247 141 251
rect 157 249 159 254
rect 164 249 166 254
rect 228 258 230 263
rect 187 247 189 251
rect 215 247 217 251
rect 238 249 240 254
rect 245 249 247 254
rect 314 270 316 282
rect 324 280 326 291
rect 344 288 346 291
rect 357 288 359 291
rect 344 286 350 288
rect 344 284 346 286
rect 348 284 350 286
rect 344 282 350 284
rect 354 286 360 288
rect 354 284 356 286
rect 358 284 360 286
rect 354 282 360 284
rect 324 278 330 280
rect 344 279 346 282
rect 324 276 326 278
rect 328 276 330 278
rect 324 274 330 276
rect 324 270 326 274
rect 354 270 356 282
rect 364 280 366 291
rect 385 289 391 291
rect 364 278 370 280
rect 364 276 366 278
rect 368 276 370 278
rect 385 276 387 289
rect 395 285 397 298
rect 474 305 476 310
rect 391 283 397 285
rect 391 281 393 283
rect 395 281 397 283
rect 405 288 407 291
rect 415 288 417 291
rect 435 288 437 291
rect 442 288 444 291
rect 453 288 455 297
rect 487 304 489 309
rect 494 304 496 309
rect 514 305 516 310
rect 635 311 637 315
rect 646 311 648 315
rect 653 311 655 315
rect 527 304 529 309
rect 534 304 536 309
rect 554 304 556 309
rect 561 304 563 309
rect 574 305 576 310
rect 594 304 596 309
rect 601 304 603 309
rect 614 305 616 310
rect 474 288 476 291
rect 487 288 489 291
rect 405 286 411 288
rect 405 284 407 286
rect 409 284 411 286
rect 405 282 411 284
rect 415 286 437 288
rect 415 284 426 286
rect 428 284 433 286
rect 435 284 437 286
rect 415 282 437 284
rect 441 286 447 288
rect 441 284 443 286
rect 445 284 447 286
rect 441 282 447 284
rect 451 286 457 288
rect 451 284 453 286
rect 455 284 457 286
rect 451 282 457 284
rect 474 286 480 288
rect 474 284 476 286
rect 478 284 480 286
rect 474 282 480 284
rect 484 286 490 288
rect 484 284 486 286
rect 488 284 490 286
rect 484 282 490 284
rect 391 279 400 281
rect 408 279 410 282
rect 415 279 417 282
rect 433 279 435 282
rect 443 279 445 282
rect 453 279 455 282
rect 474 279 476 282
rect 398 276 400 279
rect 364 274 370 276
rect 364 270 366 274
rect 398 258 400 263
rect 263 247 265 251
rect 273 247 275 251
rect 283 247 285 251
rect 304 247 306 251
rect 314 247 316 251
rect 324 247 326 251
rect 344 247 346 251
rect 354 247 356 251
rect 364 247 366 251
rect 385 247 387 251
rect 408 249 410 254
rect 415 249 417 254
rect 484 270 486 282
rect 494 280 496 291
rect 514 288 516 291
rect 527 288 529 291
rect 514 286 520 288
rect 514 284 516 286
rect 518 284 520 286
rect 514 282 520 284
rect 524 286 530 288
rect 524 284 526 286
rect 528 284 530 286
rect 524 282 530 284
rect 494 278 500 280
rect 514 279 516 282
rect 494 276 496 278
rect 498 276 500 278
rect 494 274 500 276
rect 494 270 496 274
rect 524 270 526 282
rect 534 280 536 291
rect 554 280 556 291
rect 561 288 563 291
rect 574 288 576 291
rect 560 286 566 288
rect 560 284 562 286
rect 564 284 566 286
rect 560 282 566 284
rect 570 286 576 288
rect 570 284 572 286
rect 574 284 576 286
rect 570 282 576 284
rect 534 278 540 280
rect 534 276 536 278
rect 538 276 540 278
rect 534 274 540 276
rect 550 278 556 280
rect 550 276 552 278
rect 554 276 556 278
rect 550 274 556 276
rect 534 270 536 274
rect 554 270 556 274
rect 564 270 566 282
rect 574 279 576 282
rect 594 280 596 291
rect 601 288 603 291
rect 614 288 616 291
rect 635 288 637 297
rect 673 305 675 310
rect 683 305 685 310
rect 693 308 695 313
rect 703 311 705 315
rect 646 288 648 291
rect 653 288 655 291
rect 673 288 675 291
rect 683 288 685 291
rect 600 286 606 288
rect 600 284 602 286
rect 604 284 606 286
rect 600 282 606 284
rect 610 286 616 288
rect 610 284 612 286
rect 614 284 616 286
rect 610 282 616 284
rect 633 286 639 288
rect 633 284 635 286
rect 637 284 639 286
rect 633 282 639 284
rect 643 286 649 288
rect 643 284 645 286
rect 647 284 649 286
rect 643 282 649 284
rect 653 286 675 288
rect 653 284 655 286
rect 657 284 662 286
rect 664 284 675 286
rect 653 282 675 284
rect 679 286 685 288
rect 679 284 681 286
rect 683 284 685 286
rect 679 282 685 284
rect 693 285 695 298
rect 703 295 705 298
rect 699 293 705 295
rect 699 291 701 293
rect 703 291 705 293
rect 699 289 705 291
rect 693 283 699 285
rect 590 278 596 280
rect 590 276 592 278
rect 594 276 596 278
rect 590 274 596 276
rect 594 270 596 274
rect 604 270 606 282
rect 614 279 616 282
rect 635 279 637 282
rect 645 279 647 282
rect 655 279 657 282
rect 673 279 675 282
rect 680 279 682 282
rect 693 281 695 283
rect 697 281 699 283
rect 690 279 699 281
rect 690 276 692 279
rect 703 276 705 289
rect 690 258 692 263
rect 433 247 435 251
rect 443 247 445 251
rect 453 247 455 251
rect 474 247 476 251
rect 484 247 486 251
rect 494 247 496 251
rect 514 247 516 251
rect 524 247 526 251
rect 534 247 536 251
rect 554 247 556 251
rect 564 247 566 251
rect 574 247 576 251
rect 594 247 596 251
rect 604 247 606 251
rect 614 247 616 251
rect 635 247 637 251
rect 645 247 647 251
rect 655 247 657 251
rect 673 249 675 254
rect 680 249 682 254
rect 703 247 705 251
rect 38 239 40 243
rect 51 239 53 243
rect 58 239 60 243
rect 79 239 81 243
rect 89 239 91 243
rect 99 239 101 243
rect 117 236 119 241
rect 124 236 126 241
rect 147 239 149 243
rect 180 239 182 243
rect 190 239 192 243
rect 200 239 202 243
rect 134 227 136 232
rect 134 211 136 214
rect 38 208 40 211
rect 51 208 53 211
rect 58 208 60 211
rect 79 208 81 211
rect 89 208 91 211
rect 99 208 101 211
rect 117 208 119 211
rect 124 208 126 211
rect 134 209 143 211
rect 38 206 44 208
rect 38 204 40 206
rect 42 204 44 206
rect 38 202 44 204
rect 48 206 54 208
rect 48 204 50 206
rect 52 204 54 206
rect 48 202 54 204
rect 58 206 67 208
rect 58 204 63 206
rect 65 204 67 206
rect 58 202 67 204
rect 77 206 83 208
rect 77 204 79 206
rect 81 204 83 206
rect 77 202 83 204
rect 87 206 93 208
rect 87 204 89 206
rect 91 204 93 206
rect 87 202 93 204
rect 97 206 119 208
rect 97 204 99 206
rect 101 204 106 206
rect 108 204 119 206
rect 97 202 119 204
rect 123 206 129 208
rect 123 204 125 206
rect 127 204 129 206
rect 123 202 129 204
rect 38 199 40 202
rect 48 194 50 202
rect 58 196 60 202
rect 79 193 81 202
rect 90 199 92 202
rect 97 199 99 202
rect 117 199 119 202
rect 127 199 129 202
rect 137 207 139 209
rect 141 207 143 209
rect 137 205 143 207
rect 38 180 40 185
rect 48 181 50 186
rect 58 184 60 188
rect 137 192 139 205
rect 147 201 149 214
rect 218 236 220 241
rect 225 236 227 241
rect 248 239 250 243
rect 282 239 284 243
rect 292 239 294 243
rect 302 239 304 243
rect 235 227 237 232
rect 235 211 237 214
rect 180 208 182 211
rect 190 208 192 211
rect 200 208 202 211
rect 218 208 220 211
rect 225 208 227 211
rect 235 209 244 211
rect 178 206 184 208
rect 178 204 180 206
rect 182 204 184 206
rect 178 202 184 204
rect 188 206 194 208
rect 188 204 190 206
rect 192 204 194 206
rect 188 202 194 204
rect 198 206 220 208
rect 198 204 200 206
rect 202 204 207 206
rect 209 204 220 206
rect 198 202 220 204
rect 224 206 230 208
rect 224 204 226 206
rect 228 204 230 206
rect 224 202 230 204
rect 143 199 149 201
rect 143 197 145 199
rect 147 197 149 199
rect 143 195 149 197
rect 147 192 149 195
rect 180 193 182 202
rect 191 199 193 202
rect 198 199 200 202
rect 218 199 220 202
rect 228 199 230 202
rect 238 207 240 209
rect 242 207 244 209
rect 238 205 244 207
rect 117 180 119 185
rect 127 180 129 185
rect 79 175 81 179
rect 90 175 92 179
rect 97 175 99 179
rect 137 177 139 182
rect 238 192 240 205
rect 248 201 250 214
rect 320 236 322 241
rect 327 236 329 241
rect 350 239 352 243
rect 382 239 384 243
rect 337 227 339 232
rect 337 211 339 214
rect 282 208 284 211
rect 292 208 294 211
rect 302 208 304 211
rect 320 208 322 211
rect 327 208 329 211
rect 337 209 346 211
rect 280 206 286 208
rect 280 204 282 206
rect 284 204 286 206
rect 280 202 286 204
rect 290 206 296 208
rect 290 204 292 206
rect 294 204 296 206
rect 290 202 296 204
rect 300 206 322 208
rect 300 204 302 206
rect 304 204 309 206
rect 311 204 322 206
rect 300 202 322 204
rect 326 206 332 208
rect 326 204 328 206
rect 330 204 332 206
rect 326 202 332 204
rect 244 199 250 201
rect 244 197 246 199
rect 248 197 250 199
rect 244 195 250 197
rect 248 192 250 195
rect 282 193 284 202
rect 293 199 295 202
rect 300 199 302 202
rect 320 199 322 202
rect 330 199 332 202
rect 340 207 342 209
rect 344 207 346 209
rect 340 205 346 207
rect 218 180 220 185
rect 228 180 230 185
rect 147 175 149 179
rect 180 175 182 179
rect 191 175 193 179
rect 198 175 200 179
rect 238 177 240 182
rect 340 192 342 205
rect 350 201 352 214
rect 395 239 397 243
rect 402 239 404 243
rect 435 239 437 243
rect 445 239 447 243
rect 455 239 457 243
rect 473 236 475 241
rect 480 236 482 241
rect 503 239 505 243
rect 536 239 538 243
rect 546 239 548 243
rect 556 239 558 243
rect 490 227 492 232
rect 490 211 492 214
rect 346 199 352 201
rect 382 208 384 211
rect 395 208 397 211
rect 402 208 404 211
rect 435 208 437 211
rect 445 208 447 211
rect 455 208 457 211
rect 473 208 475 211
rect 480 208 482 211
rect 490 209 499 211
rect 382 206 388 208
rect 382 204 384 206
rect 386 204 388 206
rect 382 202 388 204
rect 392 206 398 208
rect 392 204 394 206
rect 396 204 398 206
rect 392 202 398 204
rect 402 206 411 208
rect 402 204 407 206
rect 409 204 411 206
rect 402 202 411 204
rect 433 206 439 208
rect 433 204 435 206
rect 437 204 439 206
rect 433 202 439 204
rect 443 206 449 208
rect 443 204 445 206
rect 447 204 449 206
rect 443 202 449 204
rect 453 206 475 208
rect 453 204 455 206
rect 457 204 462 206
rect 464 204 475 206
rect 453 202 475 204
rect 479 206 485 208
rect 479 204 481 206
rect 483 204 485 206
rect 479 202 485 204
rect 382 199 384 202
rect 346 197 348 199
rect 350 197 352 199
rect 346 195 352 197
rect 350 192 352 195
rect 320 180 322 185
rect 330 180 332 185
rect 248 175 250 179
rect 282 175 284 179
rect 293 175 295 179
rect 300 175 302 179
rect 340 177 342 182
rect 392 194 394 202
rect 402 196 404 202
rect 435 193 437 202
rect 446 199 448 202
rect 453 199 455 202
rect 473 199 475 202
rect 483 199 485 202
rect 493 207 495 209
rect 497 207 499 209
rect 493 205 499 207
rect 382 180 384 185
rect 392 181 394 186
rect 402 184 404 188
rect 350 175 352 179
rect 493 192 495 205
rect 503 201 505 214
rect 574 236 576 241
rect 581 236 583 241
rect 604 239 606 243
rect 635 239 637 243
rect 645 239 647 243
rect 655 239 657 243
rect 591 227 593 232
rect 591 211 593 214
rect 536 208 538 211
rect 546 208 548 211
rect 556 208 558 211
rect 574 208 576 211
rect 581 208 583 211
rect 591 209 600 211
rect 534 206 540 208
rect 534 204 536 206
rect 538 204 540 206
rect 534 202 540 204
rect 544 206 550 208
rect 544 204 546 206
rect 548 204 550 206
rect 544 202 550 204
rect 554 206 576 208
rect 554 204 556 206
rect 558 204 563 206
rect 565 204 576 206
rect 554 202 576 204
rect 580 206 586 208
rect 580 204 582 206
rect 584 204 586 206
rect 580 202 586 204
rect 499 199 505 201
rect 499 197 501 199
rect 503 197 505 199
rect 499 195 505 197
rect 503 192 505 195
rect 536 193 538 202
rect 547 199 549 202
rect 554 199 556 202
rect 574 199 576 202
rect 584 199 586 202
rect 594 207 596 209
rect 598 207 600 209
rect 594 205 600 207
rect 473 180 475 185
rect 483 180 485 185
rect 435 175 437 179
rect 446 175 448 179
rect 453 175 455 179
rect 493 177 495 182
rect 594 192 596 205
rect 604 201 606 214
rect 673 236 675 241
rect 680 236 682 241
rect 703 239 705 243
rect 690 227 692 232
rect 690 211 692 214
rect 635 208 637 211
rect 645 208 647 211
rect 655 208 657 211
rect 673 208 675 211
rect 680 208 682 211
rect 690 209 699 211
rect 633 206 639 208
rect 633 204 635 206
rect 637 204 639 206
rect 633 202 639 204
rect 643 206 649 208
rect 643 204 645 206
rect 647 204 649 206
rect 643 202 649 204
rect 653 206 675 208
rect 653 204 655 206
rect 657 204 662 206
rect 664 204 675 206
rect 653 202 675 204
rect 679 206 685 208
rect 679 204 681 206
rect 683 204 685 206
rect 679 202 685 204
rect 600 199 606 201
rect 600 197 602 199
rect 604 197 606 199
rect 600 195 606 197
rect 604 192 606 195
rect 635 193 637 202
rect 646 199 648 202
rect 653 199 655 202
rect 673 199 675 202
rect 683 199 685 202
rect 693 207 695 209
rect 697 207 699 209
rect 693 205 699 207
rect 574 180 576 185
rect 584 180 586 185
rect 503 175 505 179
rect 536 175 538 179
rect 547 175 549 179
rect 554 175 556 179
rect 594 177 596 182
rect 693 192 695 205
rect 703 201 705 214
rect 699 199 705 201
rect 699 197 701 199
rect 703 197 705 199
rect 699 195 705 197
rect 703 192 705 195
rect 673 180 675 185
rect 683 180 685 185
rect 604 175 606 179
rect 635 175 637 179
rect 646 175 648 179
rect 653 175 655 179
rect 693 177 695 182
rect 703 175 705 179
rect 40 167 42 171
rect 51 167 53 171
rect 58 167 60 171
rect 40 144 42 153
rect 78 161 80 166
rect 88 161 90 166
rect 98 164 100 169
rect 108 167 110 171
rect 181 167 183 171
rect 192 167 194 171
rect 199 167 201 171
rect 128 161 130 166
rect 51 144 53 147
rect 58 144 60 147
rect 78 144 80 147
rect 88 144 90 147
rect 38 142 44 144
rect 38 140 40 142
rect 42 140 44 142
rect 38 138 44 140
rect 48 142 54 144
rect 48 140 50 142
rect 52 140 54 142
rect 48 138 54 140
rect 58 142 80 144
rect 58 140 60 142
rect 62 140 67 142
rect 69 140 80 142
rect 58 138 80 140
rect 84 142 90 144
rect 84 140 86 142
rect 88 140 90 142
rect 84 138 90 140
rect 98 141 100 154
rect 108 151 110 154
rect 104 149 110 151
rect 104 147 106 149
rect 108 147 110 149
rect 138 160 140 165
rect 148 158 150 162
rect 104 145 110 147
rect 98 139 104 141
rect 40 135 42 138
rect 50 135 52 138
rect 60 135 62 138
rect 78 135 80 138
rect 85 135 87 138
rect 98 137 100 139
rect 102 137 104 139
rect 95 135 104 137
rect 95 132 97 135
rect 108 132 110 145
rect 128 144 130 147
rect 138 144 140 152
rect 148 144 150 150
rect 181 144 183 153
rect 219 161 221 166
rect 229 161 231 166
rect 239 164 241 169
rect 249 167 251 171
rect 281 167 283 171
rect 291 164 293 169
rect 331 167 333 171
rect 338 167 340 171
rect 349 167 351 171
rect 301 161 303 166
rect 311 161 313 166
rect 192 144 194 147
rect 199 144 201 147
rect 219 144 221 147
rect 229 144 231 147
rect 128 142 134 144
rect 128 140 130 142
rect 132 140 134 142
rect 128 138 134 140
rect 138 142 144 144
rect 138 140 140 142
rect 142 140 144 142
rect 138 138 144 140
rect 148 142 157 144
rect 148 140 153 142
rect 155 140 157 142
rect 148 138 157 140
rect 179 142 185 144
rect 179 140 181 142
rect 183 140 185 142
rect 179 138 185 140
rect 189 142 195 144
rect 189 140 191 142
rect 193 140 195 142
rect 189 138 195 140
rect 199 142 221 144
rect 199 140 201 142
rect 203 140 208 142
rect 210 140 221 142
rect 199 138 221 140
rect 225 142 231 144
rect 225 140 227 142
rect 229 140 231 142
rect 225 138 231 140
rect 239 141 241 154
rect 249 151 251 154
rect 245 149 251 151
rect 245 147 247 149
rect 249 147 251 149
rect 245 145 251 147
rect 239 139 245 141
rect 128 135 130 138
rect 141 135 143 138
rect 148 135 150 138
rect 181 135 183 138
rect 191 135 193 138
rect 201 135 203 138
rect 219 135 221 138
rect 226 135 228 138
rect 239 137 241 139
rect 243 137 245 139
rect 236 135 245 137
rect 95 114 97 119
rect 40 103 42 107
rect 50 103 52 107
rect 60 103 62 107
rect 78 105 80 110
rect 85 105 87 110
rect 108 103 110 107
rect 128 103 130 107
rect 236 132 238 135
rect 249 132 251 145
rect 281 151 283 154
rect 281 149 287 151
rect 281 147 283 149
rect 285 147 287 149
rect 281 145 287 147
rect 281 132 283 145
rect 291 141 293 154
rect 435 167 437 171
rect 446 167 448 171
rect 453 167 455 171
rect 382 161 384 166
rect 287 139 293 141
rect 287 137 289 139
rect 291 137 293 139
rect 301 144 303 147
rect 311 144 313 147
rect 331 144 333 147
rect 338 144 340 147
rect 349 144 351 153
rect 392 160 394 165
rect 402 158 404 162
rect 382 144 384 147
rect 392 144 394 152
rect 402 144 404 150
rect 435 144 437 153
rect 473 161 475 166
rect 483 161 485 166
rect 493 164 495 169
rect 503 167 505 171
rect 536 167 538 171
rect 547 167 549 171
rect 554 167 556 171
rect 446 144 448 147
rect 453 144 455 147
rect 473 144 475 147
rect 483 144 485 147
rect 301 142 307 144
rect 301 140 303 142
rect 305 140 307 142
rect 301 138 307 140
rect 311 142 333 144
rect 311 140 322 142
rect 324 140 329 142
rect 331 140 333 142
rect 311 138 333 140
rect 337 142 343 144
rect 337 140 339 142
rect 341 140 343 142
rect 337 138 343 140
rect 347 142 353 144
rect 347 140 349 142
rect 351 140 353 142
rect 347 138 353 140
rect 382 142 388 144
rect 382 140 384 142
rect 386 140 388 142
rect 382 138 388 140
rect 392 142 398 144
rect 392 140 394 142
rect 396 140 398 142
rect 392 138 398 140
rect 402 142 411 144
rect 402 140 407 142
rect 409 140 411 142
rect 402 138 411 140
rect 433 142 439 144
rect 433 140 435 142
rect 437 140 439 142
rect 433 138 439 140
rect 443 142 449 144
rect 443 140 445 142
rect 447 140 449 142
rect 443 138 449 140
rect 453 142 475 144
rect 453 140 455 142
rect 457 140 462 142
rect 464 140 475 142
rect 453 138 475 140
rect 479 142 485 144
rect 479 140 481 142
rect 483 140 485 142
rect 479 138 485 140
rect 493 141 495 154
rect 503 151 505 154
rect 499 149 505 151
rect 499 147 501 149
rect 503 147 505 149
rect 499 145 505 147
rect 493 139 499 141
rect 287 135 296 137
rect 304 135 306 138
rect 311 135 313 138
rect 329 135 331 138
rect 339 135 341 138
rect 349 135 351 138
rect 382 135 384 138
rect 395 135 397 138
rect 402 135 404 138
rect 435 135 437 138
rect 445 135 447 138
rect 455 135 457 138
rect 473 135 475 138
rect 480 135 482 138
rect 493 137 495 139
rect 497 137 499 139
rect 490 135 499 137
rect 294 132 296 135
rect 236 114 238 119
rect 141 103 143 107
rect 148 103 150 107
rect 181 103 183 107
rect 191 103 193 107
rect 201 103 203 107
rect 219 105 221 110
rect 226 105 228 110
rect 294 114 296 119
rect 249 103 251 107
rect 281 103 283 107
rect 304 105 306 110
rect 311 105 313 110
rect 329 103 331 107
rect 339 103 341 107
rect 349 103 351 107
rect 382 103 384 107
rect 490 132 492 135
rect 503 132 505 145
rect 536 144 538 153
rect 574 161 576 166
rect 584 161 586 166
rect 594 164 596 169
rect 604 167 606 171
rect 635 167 637 171
rect 646 167 648 171
rect 653 167 655 171
rect 547 144 549 147
rect 554 144 556 147
rect 574 144 576 147
rect 584 144 586 147
rect 534 142 540 144
rect 534 140 536 142
rect 538 140 540 142
rect 534 138 540 140
rect 544 142 550 144
rect 544 140 546 142
rect 548 140 550 142
rect 544 138 550 140
rect 554 142 576 144
rect 554 140 556 142
rect 558 140 563 142
rect 565 140 576 142
rect 554 138 576 140
rect 580 142 586 144
rect 580 140 582 142
rect 584 140 586 142
rect 580 138 586 140
rect 594 141 596 154
rect 604 151 606 154
rect 600 149 606 151
rect 600 147 602 149
rect 604 147 606 149
rect 600 145 606 147
rect 594 139 600 141
rect 536 135 538 138
rect 546 135 548 138
rect 556 135 558 138
rect 574 135 576 138
rect 581 135 583 138
rect 594 137 596 139
rect 598 137 600 139
rect 591 135 600 137
rect 490 114 492 119
rect 395 103 397 107
rect 402 103 404 107
rect 435 103 437 107
rect 445 103 447 107
rect 455 103 457 107
rect 473 105 475 110
rect 480 105 482 110
rect 591 132 593 135
rect 604 132 606 145
rect 635 144 637 153
rect 673 161 675 166
rect 683 161 685 166
rect 693 164 695 169
rect 703 167 705 171
rect 646 144 648 147
rect 653 144 655 147
rect 673 144 675 147
rect 683 144 685 147
rect 633 142 639 144
rect 633 140 635 142
rect 637 140 639 142
rect 633 138 639 140
rect 643 142 649 144
rect 643 140 645 142
rect 647 140 649 142
rect 643 138 649 140
rect 653 142 675 144
rect 653 140 655 142
rect 657 140 662 142
rect 664 140 675 142
rect 653 138 675 140
rect 679 142 685 144
rect 679 140 681 142
rect 683 140 685 142
rect 679 138 685 140
rect 693 141 695 154
rect 703 151 705 154
rect 699 149 705 151
rect 699 147 701 149
rect 703 147 705 149
rect 699 145 705 147
rect 693 139 699 141
rect 635 135 637 138
rect 645 135 647 138
rect 655 135 657 138
rect 673 135 675 138
rect 680 135 682 138
rect 693 137 695 139
rect 697 137 699 139
rect 690 135 699 137
rect 591 114 593 119
rect 503 103 505 107
rect 536 103 538 107
rect 546 103 548 107
rect 556 103 558 107
rect 574 105 576 110
rect 581 105 583 110
rect 690 132 692 135
rect 703 132 705 145
rect 690 114 692 119
rect 604 103 606 107
rect 635 103 637 107
rect 645 103 647 107
rect 655 103 657 107
rect 673 105 675 110
rect 680 105 682 110
rect 703 103 705 107
rect 38 95 40 99
rect 51 95 53 99
rect 58 95 60 99
rect 79 95 81 99
rect 89 95 91 99
rect 99 95 101 99
rect 117 92 119 97
rect 124 92 126 97
rect 147 95 149 99
rect 180 95 182 99
rect 190 95 192 99
rect 200 95 202 99
rect 134 83 136 88
rect 134 67 136 70
rect 38 64 40 67
rect 51 64 53 67
rect 58 64 60 67
rect 79 64 81 67
rect 89 64 91 67
rect 99 64 101 67
rect 117 64 119 67
rect 124 64 126 67
rect 134 65 143 67
rect 38 62 44 64
rect 38 60 40 62
rect 42 60 44 62
rect 38 58 44 60
rect 48 62 54 64
rect 48 60 50 62
rect 52 60 54 62
rect 48 58 54 60
rect 58 62 67 64
rect 58 60 63 62
rect 65 60 67 62
rect 58 58 67 60
rect 77 62 83 64
rect 77 60 79 62
rect 81 60 83 62
rect 77 58 83 60
rect 87 62 93 64
rect 87 60 89 62
rect 91 60 93 62
rect 87 58 93 60
rect 97 62 119 64
rect 97 60 99 62
rect 101 60 106 62
rect 108 60 119 62
rect 97 58 119 60
rect 123 62 129 64
rect 123 60 125 62
rect 127 60 129 62
rect 123 58 129 60
rect 38 55 40 58
rect 48 50 50 58
rect 58 52 60 58
rect 79 49 81 58
rect 90 55 92 58
rect 97 55 99 58
rect 117 55 119 58
rect 127 55 129 58
rect 137 63 139 65
rect 141 63 143 65
rect 137 61 143 63
rect 38 36 40 41
rect 48 37 50 42
rect 58 40 60 44
rect 137 48 139 61
rect 147 57 149 70
rect 218 92 220 97
rect 225 92 227 97
rect 248 95 250 99
rect 281 95 283 99
rect 291 95 293 99
rect 301 95 303 99
rect 235 83 237 88
rect 235 67 237 70
rect 180 64 182 67
rect 190 64 192 67
rect 200 64 202 67
rect 218 64 220 67
rect 225 64 227 67
rect 235 65 244 67
rect 178 62 184 64
rect 178 60 180 62
rect 182 60 184 62
rect 178 58 184 60
rect 188 62 194 64
rect 188 60 190 62
rect 192 60 194 62
rect 188 58 194 60
rect 198 62 220 64
rect 198 60 200 62
rect 202 60 207 62
rect 209 60 220 62
rect 198 58 220 60
rect 224 62 230 64
rect 224 60 226 62
rect 228 60 230 62
rect 224 58 230 60
rect 143 55 149 57
rect 143 53 145 55
rect 147 53 149 55
rect 143 51 149 53
rect 147 48 149 51
rect 180 49 182 58
rect 191 55 193 58
rect 198 55 200 58
rect 218 55 220 58
rect 228 55 230 58
rect 238 63 240 65
rect 242 63 244 65
rect 238 61 244 63
rect 117 36 119 41
rect 127 36 129 41
rect 79 31 81 35
rect 90 31 92 35
rect 97 31 99 35
rect 137 33 139 38
rect 238 48 240 61
rect 248 57 250 70
rect 319 92 321 97
rect 326 92 328 97
rect 349 95 351 99
rect 381 95 383 99
rect 336 83 338 88
rect 336 67 338 70
rect 281 64 283 67
rect 291 64 293 67
rect 301 64 303 67
rect 319 64 321 67
rect 326 64 328 67
rect 336 65 345 67
rect 279 62 285 64
rect 279 60 281 62
rect 283 60 285 62
rect 279 58 285 60
rect 289 62 295 64
rect 289 60 291 62
rect 293 60 295 62
rect 289 58 295 60
rect 299 62 321 64
rect 299 60 301 62
rect 303 60 308 62
rect 310 60 321 62
rect 299 58 321 60
rect 325 62 331 64
rect 325 60 327 62
rect 329 60 331 62
rect 325 58 331 60
rect 244 55 250 57
rect 244 53 246 55
rect 248 53 250 55
rect 244 51 250 53
rect 248 48 250 51
rect 281 49 283 58
rect 292 55 294 58
rect 299 55 301 58
rect 319 55 321 58
rect 329 55 331 58
rect 339 63 341 65
rect 343 63 345 65
rect 339 61 345 63
rect 218 36 220 41
rect 228 36 230 41
rect 147 31 149 35
rect 180 31 182 35
rect 191 31 193 35
rect 198 31 200 35
rect 238 33 240 38
rect 339 48 341 61
rect 349 57 351 70
rect 394 95 396 99
rect 401 95 403 99
rect 434 95 436 99
rect 444 95 446 99
rect 454 95 456 99
rect 472 92 474 97
rect 479 92 481 97
rect 502 95 504 99
rect 535 95 537 99
rect 545 95 547 99
rect 555 95 557 99
rect 489 83 491 88
rect 489 67 491 70
rect 345 55 351 57
rect 381 64 383 67
rect 394 64 396 67
rect 401 64 403 67
rect 434 64 436 67
rect 444 64 446 67
rect 454 64 456 67
rect 472 64 474 67
rect 479 64 481 67
rect 489 65 498 67
rect 381 62 387 64
rect 381 60 383 62
rect 385 60 387 62
rect 381 58 387 60
rect 391 62 397 64
rect 391 60 393 62
rect 395 60 397 62
rect 391 58 397 60
rect 401 62 410 64
rect 401 60 406 62
rect 408 60 410 62
rect 401 58 410 60
rect 432 62 438 64
rect 432 60 434 62
rect 436 60 438 62
rect 432 58 438 60
rect 442 62 448 64
rect 442 60 444 62
rect 446 60 448 62
rect 442 58 448 60
rect 452 62 474 64
rect 452 60 454 62
rect 456 60 461 62
rect 463 60 474 62
rect 452 58 474 60
rect 478 62 484 64
rect 478 60 480 62
rect 482 60 484 62
rect 478 58 484 60
rect 381 55 383 58
rect 345 53 347 55
rect 349 53 351 55
rect 345 51 351 53
rect 349 48 351 51
rect 319 36 321 41
rect 329 36 331 41
rect 248 31 250 35
rect 281 31 283 35
rect 292 31 294 35
rect 299 31 301 35
rect 339 33 341 38
rect 391 50 393 58
rect 401 52 403 58
rect 434 49 436 58
rect 445 55 447 58
rect 452 55 454 58
rect 472 55 474 58
rect 482 55 484 58
rect 492 63 494 65
rect 496 63 498 65
rect 492 61 498 63
rect 381 36 383 41
rect 391 37 393 42
rect 401 40 403 44
rect 349 31 351 35
rect 492 48 494 61
rect 502 57 504 70
rect 573 92 575 97
rect 580 92 582 97
rect 603 95 605 99
rect 634 95 636 99
rect 644 95 646 99
rect 654 95 656 99
rect 590 83 592 88
rect 590 67 592 70
rect 535 64 537 67
rect 545 64 547 67
rect 555 64 557 67
rect 573 64 575 67
rect 580 64 582 67
rect 590 65 599 67
rect 533 62 539 64
rect 533 60 535 62
rect 537 60 539 62
rect 533 58 539 60
rect 543 62 549 64
rect 543 60 545 62
rect 547 60 549 62
rect 543 58 549 60
rect 553 62 575 64
rect 553 60 555 62
rect 557 60 562 62
rect 564 60 575 62
rect 553 58 575 60
rect 579 62 585 64
rect 579 60 581 62
rect 583 60 585 62
rect 579 58 585 60
rect 498 55 504 57
rect 498 53 500 55
rect 502 53 504 55
rect 498 51 504 53
rect 502 48 504 51
rect 535 49 537 58
rect 546 55 548 58
rect 553 55 555 58
rect 573 55 575 58
rect 583 55 585 58
rect 593 63 595 65
rect 597 63 599 65
rect 593 61 599 63
rect 472 36 474 41
rect 482 36 484 41
rect 434 31 436 35
rect 445 31 447 35
rect 452 31 454 35
rect 492 33 494 38
rect 593 48 595 61
rect 603 57 605 70
rect 672 92 674 97
rect 679 92 681 97
rect 702 95 704 99
rect 689 83 691 88
rect 689 67 691 70
rect 634 64 636 67
rect 644 64 646 67
rect 654 64 656 67
rect 672 64 674 67
rect 679 64 681 67
rect 689 65 698 67
rect 632 62 638 64
rect 632 60 634 62
rect 636 60 638 62
rect 632 58 638 60
rect 642 62 648 64
rect 642 60 644 62
rect 646 60 648 62
rect 642 58 648 60
rect 652 62 674 64
rect 652 60 654 62
rect 656 60 661 62
rect 663 60 674 62
rect 652 58 674 60
rect 678 62 684 64
rect 678 60 680 62
rect 682 60 684 62
rect 678 58 684 60
rect 599 55 605 57
rect 599 53 601 55
rect 603 53 605 55
rect 599 51 605 53
rect 603 48 605 51
rect 634 49 636 58
rect 645 55 647 58
rect 652 55 654 58
rect 672 55 674 58
rect 682 55 684 58
rect 692 63 694 65
rect 696 63 698 65
rect 692 61 698 63
rect 573 36 575 41
rect 583 36 585 41
rect 502 31 504 35
rect 535 31 537 35
rect 546 31 548 35
rect 553 31 555 35
rect 593 33 595 38
rect 692 48 694 61
rect 702 57 704 70
rect 698 55 704 57
rect 698 53 700 55
rect 702 53 704 55
rect 698 51 704 53
rect 702 48 704 51
rect 672 36 674 41
rect 682 36 684 41
rect 603 31 605 35
rect 634 31 636 35
rect 645 31 647 35
rect 652 31 654 35
rect 692 33 694 38
rect 702 31 704 35
<< ndif >>
rect 33 336 38 343
rect 31 334 38 336
rect 31 332 33 334
rect 35 332 38 334
rect 31 330 38 332
rect 40 330 45 343
rect 47 330 58 343
rect 49 329 58 330
rect 60 341 67 343
rect 60 339 63 341
rect 65 339 67 341
rect 60 333 67 339
rect 73 336 78 343
rect 60 331 63 333
rect 65 331 67 333
rect 60 329 67 331
rect 71 334 78 336
rect 71 332 73 334
rect 75 332 78 334
rect 71 330 78 332
rect 80 330 85 343
rect 87 330 98 343
rect 49 324 56 329
rect 89 329 98 330
rect 100 341 107 343
rect 100 339 103 341
rect 105 339 107 341
rect 100 333 107 339
rect 123 337 130 343
rect 100 331 103 333
rect 105 331 107 333
rect 100 329 107 331
rect 112 334 119 337
rect 112 332 114 334
rect 116 332 119 334
rect 112 330 119 332
rect 89 324 96 329
rect 49 322 52 324
rect 54 322 56 324
rect 49 320 56 322
rect 89 322 92 324
rect 94 322 96 324
rect 114 323 119 330
rect 121 327 130 337
rect 121 325 125 327
rect 127 325 130 327
rect 121 323 130 325
rect 132 323 137 343
rect 139 336 144 343
rect 150 341 157 343
rect 150 339 152 341
rect 154 339 157 341
rect 139 334 146 336
rect 139 332 142 334
rect 144 332 146 334
rect 139 330 146 332
rect 150 334 157 339
rect 150 332 152 334
rect 154 332 157 334
rect 139 323 144 330
rect 150 329 157 332
rect 159 341 167 343
rect 159 339 162 341
rect 164 339 167 341
rect 159 329 167 339
rect 169 336 174 343
rect 230 336 235 343
rect 169 333 177 336
rect 169 331 172 333
rect 174 331 177 333
rect 169 329 177 331
rect 172 326 177 329
rect 179 330 187 336
rect 179 328 182 330
rect 184 328 187 330
rect 179 326 187 328
rect 89 320 96 322
rect 182 323 187 326
rect 189 334 196 336
rect 189 332 192 334
rect 194 332 196 334
rect 189 330 196 332
rect 208 334 215 336
rect 208 332 210 334
rect 212 332 215 334
rect 208 330 215 332
rect 189 323 194 330
rect 210 323 215 330
rect 217 330 225 336
rect 217 328 220 330
rect 222 328 225 330
rect 217 326 225 328
rect 227 333 235 336
rect 227 331 230 333
rect 232 331 235 333
rect 227 329 235 331
rect 237 341 245 343
rect 237 339 240 341
rect 242 339 245 341
rect 237 329 245 339
rect 247 341 254 343
rect 247 339 250 341
rect 252 339 254 341
rect 247 334 254 339
rect 260 336 265 343
rect 247 332 250 334
rect 252 332 254 334
rect 247 329 254 332
rect 258 334 265 336
rect 258 332 260 334
rect 262 332 265 334
rect 258 330 265 332
rect 227 326 232 329
rect 217 323 222 326
rect 260 323 265 330
rect 267 323 272 343
rect 274 337 281 343
rect 297 341 304 343
rect 297 339 299 341
rect 301 339 304 341
rect 274 327 283 337
rect 274 325 277 327
rect 279 325 283 327
rect 274 323 283 325
rect 285 334 292 337
rect 285 332 288 334
rect 290 332 292 334
rect 285 330 292 332
rect 297 333 304 339
rect 297 331 299 333
rect 301 331 304 333
rect 285 323 290 330
rect 297 329 304 331
rect 306 330 317 343
rect 319 330 324 343
rect 326 336 331 343
rect 337 341 344 343
rect 337 339 339 341
rect 341 339 344 341
rect 326 334 333 336
rect 326 332 329 334
rect 331 332 333 334
rect 326 330 333 332
rect 337 333 344 339
rect 337 331 339 333
rect 341 331 344 333
rect 306 329 315 330
rect 308 324 315 329
rect 337 329 344 331
rect 346 330 357 343
rect 359 330 364 343
rect 366 336 371 343
rect 400 336 405 343
rect 366 334 373 336
rect 366 332 369 334
rect 371 332 373 334
rect 366 330 373 332
rect 378 334 385 336
rect 378 332 380 334
rect 382 332 385 334
rect 378 330 385 332
rect 346 329 355 330
rect 348 324 355 329
rect 308 322 310 324
rect 312 322 315 324
rect 308 320 315 322
rect 348 322 350 324
rect 352 322 355 324
rect 380 323 385 330
rect 387 330 395 336
rect 387 328 390 330
rect 392 328 395 330
rect 387 326 395 328
rect 397 333 405 336
rect 397 331 400 333
rect 402 331 405 333
rect 397 329 405 331
rect 407 341 415 343
rect 407 339 410 341
rect 412 339 415 341
rect 407 329 415 339
rect 417 341 424 343
rect 417 339 420 341
rect 422 339 424 341
rect 417 334 424 339
rect 430 336 435 343
rect 417 332 420 334
rect 422 332 424 334
rect 417 329 424 332
rect 428 334 435 336
rect 428 332 430 334
rect 432 332 435 334
rect 428 330 435 332
rect 397 326 402 329
rect 387 323 392 326
rect 348 320 355 322
rect 430 323 435 330
rect 437 323 442 343
rect 444 337 451 343
rect 467 341 474 343
rect 467 339 469 341
rect 471 339 474 341
rect 444 327 453 337
rect 444 325 447 327
rect 449 325 453 327
rect 444 323 453 325
rect 455 334 462 337
rect 455 332 458 334
rect 460 332 462 334
rect 455 330 462 332
rect 467 333 474 339
rect 467 331 469 333
rect 471 331 474 333
rect 455 323 460 330
rect 467 329 474 331
rect 476 330 487 343
rect 489 330 494 343
rect 496 336 501 343
rect 507 341 514 343
rect 507 339 509 341
rect 511 339 514 341
rect 496 334 503 336
rect 496 332 499 334
rect 501 332 503 334
rect 496 330 503 332
rect 507 333 514 339
rect 507 331 509 333
rect 511 331 514 333
rect 476 329 485 330
rect 478 324 485 329
rect 507 329 514 331
rect 516 330 527 343
rect 529 330 534 343
rect 536 336 541 343
rect 549 336 554 343
rect 536 334 543 336
rect 536 332 539 334
rect 541 332 543 334
rect 536 330 543 332
rect 547 334 554 336
rect 547 332 549 334
rect 551 332 554 334
rect 547 330 554 332
rect 556 330 561 343
rect 563 330 574 343
rect 516 329 525 330
rect 518 324 525 329
rect 565 329 574 330
rect 576 341 583 343
rect 576 339 579 341
rect 581 339 583 341
rect 576 333 583 339
rect 589 336 594 343
rect 576 331 579 333
rect 581 331 583 333
rect 576 329 583 331
rect 587 334 594 336
rect 587 332 589 334
rect 591 332 594 334
rect 587 330 594 332
rect 596 330 601 343
rect 603 330 614 343
rect 478 322 480 324
rect 482 322 485 324
rect 478 320 485 322
rect 518 322 520 324
rect 522 322 525 324
rect 518 320 525 322
rect 565 324 572 329
rect 605 329 614 330
rect 616 341 623 343
rect 616 339 619 341
rect 621 339 623 341
rect 616 333 623 339
rect 639 337 646 343
rect 616 331 619 333
rect 621 331 623 333
rect 616 329 623 331
rect 628 334 635 337
rect 628 332 630 334
rect 632 332 635 334
rect 628 330 635 332
rect 605 324 612 329
rect 565 322 568 324
rect 570 322 572 324
rect 565 320 572 322
rect 605 322 608 324
rect 610 322 612 324
rect 630 323 635 330
rect 637 327 646 337
rect 637 325 641 327
rect 643 325 646 327
rect 637 323 646 325
rect 648 323 653 343
rect 655 336 660 343
rect 666 341 673 343
rect 666 339 668 341
rect 670 339 673 341
rect 655 334 662 336
rect 655 332 658 334
rect 660 332 662 334
rect 655 330 662 332
rect 666 334 673 339
rect 666 332 668 334
rect 670 332 673 334
rect 655 323 660 330
rect 666 329 673 332
rect 675 341 683 343
rect 675 339 678 341
rect 680 339 683 341
rect 675 329 683 339
rect 685 336 690 343
rect 685 333 693 336
rect 685 331 688 333
rect 690 331 693 333
rect 685 329 693 331
rect 688 326 693 329
rect 695 330 703 336
rect 695 328 698 330
rect 700 328 703 330
rect 695 326 703 328
rect 605 320 612 322
rect 698 323 703 326
rect 705 334 712 336
rect 705 332 708 334
rect 710 332 712 334
rect 705 330 712 332
rect 705 323 710 330
rect 49 312 56 314
rect 49 310 52 312
rect 54 310 56 312
rect 89 312 96 314
rect 89 310 92 312
rect 94 310 96 312
rect 49 305 56 310
rect 49 304 58 305
rect 31 302 38 304
rect 31 300 33 302
rect 35 300 38 302
rect 31 298 38 300
rect 33 291 38 298
rect 40 291 45 304
rect 47 291 58 304
rect 60 303 67 305
rect 89 305 96 310
rect 89 304 98 305
rect 60 301 63 303
rect 65 301 67 303
rect 60 295 67 301
rect 71 302 78 304
rect 71 300 73 302
rect 75 300 78 302
rect 71 298 78 300
rect 60 293 63 295
rect 65 293 67 295
rect 60 291 67 293
rect 73 291 78 298
rect 80 291 85 304
rect 87 291 98 304
rect 100 303 107 305
rect 114 304 119 311
rect 100 301 103 303
rect 105 301 107 303
rect 100 295 107 301
rect 112 302 119 304
rect 112 300 114 302
rect 116 300 119 302
rect 112 297 119 300
rect 121 309 130 311
rect 121 307 125 309
rect 127 307 130 309
rect 121 297 130 307
rect 100 293 103 295
rect 105 293 107 295
rect 100 291 107 293
rect 123 291 130 297
rect 132 291 137 311
rect 139 304 144 311
rect 182 308 187 311
rect 172 305 177 308
rect 139 302 146 304
rect 139 300 142 302
rect 144 300 146 302
rect 139 298 146 300
rect 150 302 157 305
rect 150 300 152 302
rect 154 300 157 302
rect 139 291 144 298
rect 150 295 157 300
rect 150 293 152 295
rect 154 293 157 295
rect 150 291 157 293
rect 159 295 167 305
rect 159 293 162 295
rect 164 293 167 295
rect 159 291 167 293
rect 169 303 177 305
rect 169 301 172 303
rect 174 301 177 303
rect 169 298 177 301
rect 179 306 187 308
rect 179 304 182 306
rect 184 304 187 306
rect 179 298 187 304
rect 189 304 194 311
rect 210 304 215 311
rect 189 302 196 304
rect 189 300 192 302
rect 194 300 196 302
rect 189 298 196 300
rect 208 302 215 304
rect 208 300 210 302
rect 212 300 215 302
rect 208 298 215 300
rect 217 308 222 311
rect 308 312 315 314
rect 217 306 225 308
rect 217 304 220 306
rect 222 304 225 306
rect 217 298 225 304
rect 227 305 232 308
rect 227 303 235 305
rect 227 301 230 303
rect 232 301 235 303
rect 227 298 235 301
rect 169 291 174 298
rect 230 291 235 298
rect 237 295 245 305
rect 237 293 240 295
rect 242 293 245 295
rect 237 291 245 293
rect 247 302 254 305
rect 260 304 265 311
rect 247 300 250 302
rect 252 300 254 302
rect 247 295 254 300
rect 258 302 265 304
rect 258 300 260 302
rect 262 300 265 302
rect 258 298 265 300
rect 247 293 250 295
rect 252 293 254 295
rect 247 291 254 293
rect 260 291 265 298
rect 267 291 272 311
rect 274 309 283 311
rect 274 307 277 309
rect 279 307 283 309
rect 274 297 283 307
rect 285 304 290 311
rect 308 310 310 312
rect 312 310 315 312
rect 348 312 355 314
rect 348 310 350 312
rect 352 310 355 312
rect 308 305 315 310
rect 285 302 292 304
rect 285 300 288 302
rect 290 300 292 302
rect 285 297 292 300
rect 297 303 304 305
rect 297 301 299 303
rect 301 301 304 303
rect 274 291 281 297
rect 297 295 304 301
rect 297 293 299 295
rect 301 293 304 295
rect 297 291 304 293
rect 306 304 315 305
rect 348 305 355 310
rect 306 291 317 304
rect 319 291 324 304
rect 326 302 333 304
rect 326 300 329 302
rect 331 300 333 302
rect 326 298 333 300
rect 337 303 344 305
rect 337 301 339 303
rect 341 301 344 303
rect 326 291 331 298
rect 337 295 344 301
rect 337 293 339 295
rect 341 293 344 295
rect 337 291 344 293
rect 346 304 355 305
rect 380 304 385 311
rect 346 291 357 304
rect 359 291 364 304
rect 366 302 373 304
rect 366 300 369 302
rect 371 300 373 302
rect 366 298 373 300
rect 378 302 385 304
rect 378 300 380 302
rect 382 300 385 302
rect 378 298 385 300
rect 387 308 392 311
rect 478 312 485 314
rect 387 306 395 308
rect 387 304 390 306
rect 392 304 395 306
rect 387 298 395 304
rect 397 305 402 308
rect 397 303 405 305
rect 397 301 400 303
rect 402 301 405 303
rect 397 298 405 301
rect 366 291 371 298
rect 400 291 405 298
rect 407 295 415 305
rect 407 293 410 295
rect 412 293 415 295
rect 407 291 415 293
rect 417 302 424 305
rect 430 304 435 311
rect 417 300 420 302
rect 422 300 424 302
rect 417 295 424 300
rect 428 302 435 304
rect 428 300 430 302
rect 432 300 435 302
rect 428 298 435 300
rect 417 293 420 295
rect 422 293 424 295
rect 417 291 424 293
rect 430 291 435 298
rect 437 291 442 311
rect 444 309 453 311
rect 444 307 447 309
rect 449 307 453 309
rect 444 297 453 307
rect 455 304 460 311
rect 478 310 480 312
rect 482 310 485 312
rect 518 312 525 314
rect 518 310 520 312
rect 522 310 525 312
rect 478 305 485 310
rect 455 302 462 304
rect 455 300 458 302
rect 460 300 462 302
rect 455 297 462 300
rect 467 303 474 305
rect 467 301 469 303
rect 471 301 474 303
rect 444 291 451 297
rect 467 295 474 301
rect 467 293 469 295
rect 471 293 474 295
rect 467 291 474 293
rect 476 304 485 305
rect 518 305 525 310
rect 565 312 572 314
rect 565 310 568 312
rect 570 310 572 312
rect 605 312 612 314
rect 605 310 608 312
rect 610 310 612 312
rect 476 291 487 304
rect 489 291 494 304
rect 496 302 503 304
rect 496 300 499 302
rect 501 300 503 302
rect 496 298 503 300
rect 507 303 514 305
rect 507 301 509 303
rect 511 301 514 303
rect 496 291 501 298
rect 507 295 514 301
rect 507 293 509 295
rect 511 293 514 295
rect 507 291 514 293
rect 516 304 525 305
rect 565 305 572 310
rect 565 304 574 305
rect 516 291 527 304
rect 529 291 534 304
rect 536 302 543 304
rect 536 300 539 302
rect 541 300 543 302
rect 536 298 543 300
rect 547 302 554 304
rect 547 300 549 302
rect 551 300 554 302
rect 547 298 554 300
rect 536 291 541 298
rect 549 291 554 298
rect 556 291 561 304
rect 563 291 574 304
rect 576 303 583 305
rect 605 305 612 310
rect 605 304 614 305
rect 576 301 579 303
rect 581 301 583 303
rect 576 295 583 301
rect 587 302 594 304
rect 587 300 589 302
rect 591 300 594 302
rect 587 298 594 300
rect 576 293 579 295
rect 581 293 583 295
rect 576 291 583 293
rect 589 291 594 298
rect 596 291 601 304
rect 603 291 614 304
rect 616 303 623 305
rect 630 304 635 311
rect 616 301 619 303
rect 621 301 623 303
rect 616 295 623 301
rect 628 302 635 304
rect 628 300 630 302
rect 632 300 635 302
rect 628 297 635 300
rect 637 309 646 311
rect 637 307 641 309
rect 643 307 646 309
rect 637 297 646 307
rect 616 293 619 295
rect 621 293 623 295
rect 616 291 623 293
rect 639 291 646 297
rect 648 291 653 311
rect 655 304 660 311
rect 698 308 703 311
rect 688 305 693 308
rect 655 302 662 304
rect 655 300 658 302
rect 660 300 662 302
rect 655 298 662 300
rect 666 302 673 305
rect 666 300 668 302
rect 670 300 673 302
rect 655 291 660 298
rect 666 295 673 300
rect 666 293 668 295
rect 670 293 673 295
rect 666 291 673 293
rect 675 295 683 305
rect 675 293 678 295
rect 680 293 683 295
rect 675 291 683 293
rect 685 303 693 305
rect 685 301 688 303
rect 690 301 693 303
rect 685 298 693 301
rect 695 306 703 308
rect 695 304 698 306
rect 700 304 703 306
rect 695 298 703 304
rect 705 304 710 311
rect 705 302 712 304
rect 705 300 708 302
rect 710 300 712 302
rect 705 298 712 300
rect 685 291 690 298
rect 31 197 38 199
rect 31 195 33 197
rect 35 195 38 197
rect 31 190 38 195
rect 31 188 33 190
rect 35 188 38 190
rect 31 185 38 188
rect 40 194 45 199
rect 53 194 58 196
rect 40 190 48 194
rect 40 188 43 190
rect 45 188 48 190
rect 40 186 48 188
rect 50 192 58 194
rect 50 190 53 192
rect 55 190 58 192
rect 50 188 58 190
rect 60 192 67 196
rect 83 193 90 199
rect 60 190 63 192
rect 65 190 67 192
rect 60 188 67 190
rect 72 190 79 193
rect 72 188 74 190
rect 76 188 79 190
rect 50 186 55 188
rect 40 185 45 186
rect 72 186 79 188
rect 74 179 79 186
rect 81 183 90 193
rect 81 181 85 183
rect 87 181 90 183
rect 81 179 90 181
rect 92 179 97 199
rect 99 192 104 199
rect 110 197 117 199
rect 110 195 112 197
rect 114 195 117 197
rect 99 190 106 192
rect 99 188 102 190
rect 104 188 106 190
rect 99 186 106 188
rect 110 190 117 195
rect 110 188 112 190
rect 114 188 117 190
rect 99 179 104 186
rect 110 185 117 188
rect 119 197 127 199
rect 119 195 122 197
rect 124 195 127 197
rect 119 185 127 195
rect 129 192 134 199
rect 184 193 191 199
rect 129 189 137 192
rect 129 187 132 189
rect 134 187 137 189
rect 129 185 137 187
rect 132 182 137 185
rect 139 186 147 192
rect 139 184 142 186
rect 144 184 147 186
rect 139 182 147 184
rect 142 179 147 182
rect 149 190 156 192
rect 149 188 152 190
rect 154 188 156 190
rect 149 186 156 188
rect 173 190 180 193
rect 173 188 175 190
rect 177 188 180 190
rect 173 186 180 188
rect 149 179 154 186
rect 175 179 180 186
rect 182 183 191 193
rect 182 181 186 183
rect 188 181 191 183
rect 182 179 191 181
rect 193 179 198 199
rect 200 192 205 199
rect 211 197 218 199
rect 211 195 213 197
rect 215 195 218 197
rect 200 190 207 192
rect 200 188 203 190
rect 205 188 207 190
rect 200 186 207 188
rect 211 190 218 195
rect 211 188 213 190
rect 215 188 218 190
rect 200 179 205 186
rect 211 185 218 188
rect 220 197 228 199
rect 220 195 223 197
rect 225 195 228 197
rect 220 185 228 195
rect 230 192 235 199
rect 286 193 293 199
rect 230 189 238 192
rect 230 187 233 189
rect 235 187 238 189
rect 230 185 238 187
rect 233 182 238 185
rect 240 186 248 192
rect 240 184 243 186
rect 245 184 248 186
rect 240 182 248 184
rect 243 179 248 182
rect 250 190 257 192
rect 250 188 253 190
rect 255 188 257 190
rect 250 186 257 188
rect 275 190 282 193
rect 275 188 277 190
rect 279 188 282 190
rect 275 186 282 188
rect 250 179 255 186
rect 277 179 282 186
rect 284 183 293 193
rect 284 181 288 183
rect 290 181 293 183
rect 284 179 293 181
rect 295 179 300 199
rect 302 192 307 199
rect 313 197 320 199
rect 313 195 315 197
rect 317 195 320 197
rect 302 190 309 192
rect 302 188 305 190
rect 307 188 309 190
rect 302 186 309 188
rect 313 190 320 195
rect 313 188 315 190
rect 317 188 320 190
rect 302 179 307 186
rect 313 185 320 188
rect 322 197 330 199
rect 322 195 325 197
rect 327 195 330 197
rect 322 185 330 195
rect 332 192 337 199
rect 375 197 382 199
rect 375 195 377 197
rect 379 195 382 197
rect 332 189 340 192
rect 332 187 335 189
rect 337 187 340 189
rect 332 185 340 187
rect 335 182 340 185
rect 342 186 350 192
rect 342 184 345 186
rect 347 184 350 186
rect 342 182 350 184
rect 345 179 350 182
rect 352 190 359 192
rect 352 188 355 190
rect 357 188 359 190
rect 352 186 359 188
rect 375 190 382 195
rect 375 188 377 190
rect 379 188 382 190
rect 352 179 357 186
rect 375 185 382 188
rect 384 194 389 199
rect 397 194 402 196
rect 384 190 392 194
rect 384 188 387 190
rect 389 188 392 190
rect 384 186 392 188
rect 394 192 402 194
rect 394 190 397 192
rect 399 190 402 192
rect 394 188 402 190
rect 404 192 411 196
rect 439 193 446 199
rect 404 190 407 192
rect 409 190 411 192
rect 404 188 411 190
rect 428 190 435 193
rect 428 188 430 190
rect 432 188 435 190
rect 394 186 399 188
rect 384 185 389 186
rect 428 186 435 188
rect 430 179 435 186
rect 437 183 446 193
rect 437 181 441 183
rect 443 181 446 183
rect 437 179 446 181
rect 448 179 453 199
rect 455 192 460 199
rect 466 197 473 199
rect 466 195 468 197
rect 470 195 473 197
rect 455 190 462 192
rect 455 188 458 190
rect 460 188 462 190
rect 455 186 462 188
rect 466 190 473 195
rect 466 188 468 190
rect 470 188 473 190
rect 455 179 460 186
rect 466 185 473 188
rect 475 197 483 199
rect 475 195 478 197
rect 480 195 483 197
rect 475 185 483 195
rect 485 192 490 199
rect 540 193 547 199
rect 485 189 493 192
rect 485 187 488 189
rect 490 187 493 189
rect 485 185 493 187
rect 488 182 493 185
rect 495 186 503 192
rect 495 184 498 186
rect 500 184 503 186
rect 495 182 503 184
rect 498 179 503 182
rect 505 190 512 192
rect 505 188 508 190
rect 510 188 512 190
rect 505 186 512 188
rect 529 190 536 193
rect 529 188 531 190
rect 533 188 536 190
rect 529 186 536 188
rect 505 179 510 186
rect 531 179 536 186
rect 538 183 547 193
rect 538 181 542 183
rect 544 181 547 183
rect 538 179 547 181
rect 549 179 554 199
rect 556 192 561 199
rect 567 197 574 199
rect 567 195 569 197
rect 571 195 574 197
rect 556 190 563 192
rect 556 188 559 190
rect 561 188 563 190
rect 556 186 563 188
rect 567 190 574 195
rect 567 188 569 190
rect 571 188 574 190
rect 556 179 561 186
rect 567 185 574 188
rect 576 197 584 199
rect 576 195 579 197
rect 581 195 584 197
rect 576 185 584 195
rect 586 192 591 199
rect 639 193 646 199
rect 586 189 594 192
rect 586 187 589 189
rect 591 187 594 189
rect 586 185 594 187
rect 589 182 594 185
rect 596 186 604 192
rect 596 184 599 186
rect 601 184 604 186
rect 596 182 604 184
rect 599 179 604 182
rect 606 190 613 192
rect 606 188 609 190
rect 611 188 613 190
rect 606 186 613 188
rect 628 190 635 193
rect 628 188 630 190
rect 632 188 635 190
rect 628 186 635 188
rect 606 179 611 186
rect 630 179 635 186
rect 637 183 646 193
rect 637 181 641 183
rect 643 181 646 183
rect 637 179 646 181
rect 648 179 653 199
rect 655 192 660 199
rect 666 197 673 199
rect 666 195 668 197
rect 670 195 673 197
rect 655 190 662 192
rect 655 188 658 190
rect 660 188 662 190
rect 655 186 662 188
rect 666 190 673 195
rect 666 188 668 190
rect 670 188 673 190
rect 655 179 660 186
rect 666 185 673 188
rect 675 197 683 199
rect 675 195 678 197
rect 680 195 683 197
rect 675 185 683 195
rect 685 192 690 199
rect 685 189 693 192
rect 685 187 688 189
rect 690 187 693 189
rect 685 185 693 187
rect 688 182 693 185
rect 695 186 703 192
rect 695 184 698 186
rect 700 184 703 186
rect 695 182 703 184
rect 698 179 703 182
rect 705 190 712 192
rect 705 188 708 190
rect 710 188 712 190
rect 705 186 712 188
rect 705 179 710 186
rect 35 160 40 167
rect 33 158 40 160
rect 33 156 35 158
rect 37 156 40 158
rect 33 153 40 156
rect 42 165 51 167
rect 42 163 46 165
rect 48 163 51 165
rect 42 153 51 163
rect 44 147 51 153
rect 53 147 58 167
rect 60 160 65 167
rect 103 164 108 167
rect 93 161 98 164
rect 60 158 67 160
rect 60 156 63 158
rect 65 156 67 158
rect 60 154 67 156
rect 71 158 78 161
rect 71 156 73 158
rect 75 156 78 158
rect 60 147 65 154
rect 71 151 78 156
rect 71 149 73 151
rect 75 149 78 151
rect 71 147 78 149
rect 80 151 88 161
rect 80 149 83 151
rect 85 149 88 151
rect 80 147 88 149
rect 90 159 98 161
rect 90 157 93 159
rect 95 157 98 159
rect 90 154 98 157
rect 100 162 108 164
rect 100 160 103 162
rect 105 160 108 162
rect 100 154 108 160
rect 110 160 115 167
rect 110 158 117 160
rect 110 156 113 158
rect 115 156 117 158
rect 110 154 117 156
rect 121 158 128 161
rect 121 156 123 158
rect 125 156 128 158
rect 90 147 95 154
rect 121 151 128 156
rect 121 149 123 151
rect 125 149 128 151
rect 121 147 128 149
rect 130 160 135 161
rect 130 158 138 160
rect 130 156 133 158
rect 135 156 138 158
rect 130 152 138 156
rect 140 158 145 160
rect 176 160 181 167
rect 174 158 181 160
rect 140 156 148 158
rect 140 154 143 156
rect 145 154 148 156
rect 140 152 148 154
rect 130 147 135 152
rect 143 150 148 152
rect 150 156 157 158
rect 150 154 153 156
rect 155 154 157 156
rect 150 150 157 154
rect 174 156 176 158
rect 178 156 181 158
rect 174 153 181 156
rect 183 165 192 167
rect 183 163 187 165
rect 189 163 192 165
rect 183 153 192 163
rect 185 147 192 153
rect 194 147 199 167
rect 201 160 206 167
rect 244 164 249 167
rect 234 161 239 164
rect 201 158 208 160
rect 201 156 204 158
rect 206 156 208 158
rect 201 154 208 156
rect 212 158 219 161
rect 212 156 214 158
rect 216 156 219 158
rect 201 147 206 154
rect 212 151 219 156
rect 212 149 214 151
rect 216 149 219 151
rect 212 147 219 149
rect 221 151 229 161
rect 221 149 224 151
rect 226 149 229 151
rect 221 147 229 149
rect 231 159 239 161
rect 231 157 234 159
rect 236 157 239 159
rect 231 154 239 157
rect 241 162 249 164
rect 241 160 244 162
rect 246 160 249 162
rect 241 154 249 160
rect 251 160 256 167
rect 276 160 281 167
rect 251 158 258 160
rect 251 156 254 158
rect 256 156 258 158
rect 251 154 258 156
rect 274 158 281 160
rect 274 156 276 158
rect 278 156 281 158
rect 274 154 281 156
rect 283 164 288 167
rect 283 162 291 164
rect 283 160 286 162
rect 288 160 291 162
rect 283 154 291 160
rect 293 161 298 164
rect 293 159 301 161
rect 293 157 296 159
rect 298 157 301 159
rect 293 154 301 157
rect 231 147 236 154
rect 296 147 301 154
rect 303 151 311 161
rect 303 149 306 151
rect 308 149 311 151
rect 303 147 311 149
rect 313 158 320 161
rect 326 160 331 167
rect 313 156 316 158
rect 318 156 320 158
rect 313 151 320 156
rect 324 158 331 160
rect 324 156 326 158
rect 328 156 331 158
rect 324 154 331 156
rect 313 149 316 151
rect 318 149 320 151
rect 313 147 320 149
rect 326 147 331 154
rect 333 147 338 167
rect 340 165 349 167
rect 340 163 343 165
rect 345 163 349 165
rect 340 153 349 163
rect 351 160 356 167
rect 351 158 358 160
rect 351 156 354 158
rect 356 156 358 158
rect 351 153 358 156
rect 375 158 382 161
rect 375 156 377 158
rect 379 156 382 158
rect 340 147 347 153
rect 375 151 382 156
rect 375 149 377 151
rect 379 149 382 151
rect 375 147 382 149
rect 384 160 389 161
rect 384 158 392 160
rect 384 156 387 158
rect 389 156 392 158
rect 384 152 392 156
rect 394 158 399 160
rect 430 160 435 167
rect 428 158 435 160
rect 394 156 402 158
rect 394 154 397 156
rect 399 154 402 156
rect 394 152 402 154
rect 384 147 389 152
rect 397 150 402 152
rect 404 156 411 158
rect 404 154 407 156
rect 409 154 411 156
rect 404 150 411 154
rect 428 156 430 158
rect 432 156 435 158
rect 428 153 435 156
rect 437 165 446 167
rect 437 163 441 165
rect 443 163 446 165
rect 437 153 446 163
rect 439 147 446 153
rect 448 147 453 167
rect 455 160 460 167
rect 498 164 503 167
rect 488 161 493 164
rect 455 158 462 160
rect 455 156 458 158
rect 460 156 462 158
rect 455 154 462 156
rect 466 158 473 161
rect 466 156 468 158
rect 470 156 473 158
rect 455 147 460 154
rect 466 151 473 156
rect 466 149 468 151
rect 470 149 473 151
rect 466 147 473 149
rect 475 151 483 161
rect 475 149 478 151
rect 480 149 483 151
rect 475 147 483 149
rect 485 159 493 161
rect 485 157 488 159
rect 490 157 493 159
rect 485 154 493 157
rect 495 162 503 164
rect 495 160 498 162
rect 500 160 503 162
rect 495 154 503 160
rect 505 160 510 167
rect 531 160 536 167
rect 505 158 512 160
rect 505 156 508 158
rect 510 156 512 158
rect 505 154 512 156
rect 529 158 536 160
rect 529 156 531 158
rect 533 156 536 158
rect 485 147 490 154
rect 529 153 536 156
rect 538 165 547 167
rect 538 163 542 165
rect 544 163 547 165
rect 538 153 547 163
rect 540 147 547 153
rect 549 147 554 167
rect 556 160 561 167
rect 599 164 604 167
rect 589 161 594 164
rect 556 158 563 160
rect 556 156 559 158
rect 561 156 563 158
rect 556 154 563 156
rect 567 158 574 161
rect 567 156 569 158
rect 571 156 574 158
rect 556 147 561 154
rect 567 151 574 156
rect 567 149 569 151
rect 571 149 574 151
rect 567 147 574 149
rect 576 151 584 161
rect 576 149 579 151
rect 581 149 584 151
rect 576 147 584 149
rect 586 159 594 161
rect 586 157 589 159
rect 591 157 594 159
rect 586 154 594 157
rect 596 162 604 164
rect 596 160 599 162
rect 601 160 604 162
rect 596 154 604 160
rect 606 160 611 167
rect 630 160 635 167
rect 606 158 613 160
rect 606 156 609 158
rect 611 156 613 158
rect 606 154 613 156
rect 628 158 635 160
rect 628 156 630 158
rect 632 156 635 158
rect 586 147 591 154
rect 628 153 635 156
rect 637 165 646 167
rect 637 163 641 165
rect 643 163 646 165
rect 637 153 646 163
rect 639 147 646 153
rect 648 147 653 167
rect 655 160 660 167
rect 698 164 703 167
rect 688 161 693 164
rect 655 158 662 160
rect 655 156 658 158
rect 660 156 662 158
rect 655 154 662 156
rect 666 158 673 161
rect 666 156 668 158
rect 670 156 673 158
rect 655 147 660 154
rect 666 151 673 156
rect 666 149 668 151
rect 670 149 673 151
rect 666 147 673 149
rect 675 151 683 161
rect 675 149 678 151
rect 680 149 683 151
rect 675 147 683 149
rect 685 159 693 161
rect 685 157 688 159
rect 690 157 693 159
rect 685 154 693 157
rect 695 162 703 164
rect 695 160 698 162
rect 700 160 703 162
rect 695 154 703 160
rect 705 160 710 167
rect 705 158 712 160
rect 705 156 708 158
rect 710 156 712 158
rect 705 154 712 156
rect 685 147 690 154
rect 31 53 38 55
rect 31 51 33 53
rect 35 51 38 53
rect 31 46 38 51
rect 31 44 33 46
rect 35 44 38 46
rect 31 41 38 44
rect 40 50 45 55
rect 53 50 58 52
rect 40 46 48 50
rect 40 44 43 46
rect 45 44 48 46
rect 40 42 48 44
rect 50 48 58 50
rect 50 46 53 48
rect 55 46 58 48
rect 50 44 58 46
rect 60 48 67 52
rect 83 49 90 55
rect 60 46 63 48
rect 65 46 67 48
rect 60 44 67 46
rect 72 46 79 49
rect 72 44 74 46
rect 76 44 79 46
rect 50 42 55 44
rect 40 41 45 42
rect 72 42 79 44
rect 74 35 79 42
rect 81 39 90 49
rect 81 37 85 39
rect 87 37 90 39
rect 81 35 90 37
rect 92 35 97 55
rect 99 48 104 55
rect 110 53 117 55
rect 110 51 112 53
rect 114 51 117 53
rect 99 46 106 48
rect 99 44 102 46
rect 104 44 106 46
rect 99 42 106 44
rect 110 46 117 51
rect 110 44 112 46
rect 114 44 117 46
rect 99 35 104 42
rect 110 41 117 44
rect 119 53 127 55
rect 119 51 122 53
rect 124 51 127 53
rect 119 41 127 51
rect 129 48 134 55
rect 184 49 191 55
rect 129 45 137 48
rect 129 43 132 45
rect 134 43 137 45
rect 129 41 137 43
rect 132 38 137 41
rect 139 42 147 48
rect 139 40 142 42
rect 144 40 147 42
rect 139 38 147 40
rect 142 35 147 38
rect 149 46 156 48
rect 149 44 152 46
rect 154 44 156 46
rect 149 42 156 44
rect 173 46 180 49
rect 173 44 175 46
rect 177 44 180 46
rect 173 42 180 44
rect 149 35 154 42
rect 175 35 180 42
rect 182 39 191 49
rect 182 37 186 39
rect 188 37 191 39
rect 182 35 191 37
rect 193 35 198 55
rect 200 48 205 55
rect 211 53 218 55
rect 211 51 213 53
rect 215 51 218 53
rect 200 46 207 48
rect 200 44 203 46
rect 205 44 207 46
rect 200 42 207 44
rect 211 46 218 51
rect 211 44 213 46
rect 215 44 218 46
rect 200 35 205 42
rect 211 41 218 44
rect 220 53 228 55
rect 220 51 223 53
rect 225 51 228 53
rect 220 41 228 51
rect 230 48 235 55
rect 285 49 292 55
rect 230 45 238 48
rect 230 43 233 45
rect 235 43 238 45
rect 230 41 238 43
rect 233 38 238 41
rect 240 42 248 48
rect 240 40 243 42
rect 245 40 248 42
rect 240 38 248 40
rect 243 35 248 38
rect 250 46 257 48
rect 250 44 253 46
rect 255 44 257 46
rect 250 42 257 44
rect 274 46 281 49
rect 274 44 276 46
rect 278 44 281 46
rect 274 42 281 44
rect 250 35 255 42
rect 276 35 281 42
rect 283 39 292 49
rect 283 37 287 39
rect 289 37 292 39
rect 283 35 292 37
rect 294 35 299 55
rect 301 48 306 55
rect 312 53 319 55
rect 312 51 314 53
rect 316 51 319 53
rect 301 46 308 48
rect 301 44 304 46
rect 306 44 308 46
rect 301 42 308 44
rect 312 46 319 51
rect 312 44 314 46
rect 316 44 319 46
rect 301 35 306 42
rect 312 41 319 44
rect 321 53 329 55
rect 321 51 324 53
rect 326 51 329 53
rect 321 41 329 51
rect 331 48 336 55
rect 374 53 381 55
rect 374 51 376 53
rect 378 51 381 53
rect 331 45 339 48
rect 331 43 334 45
rect 336 43 339 45
rect 331 41 339 43
rect 334 38 339 41
rect 341 42 349 48
rect 341 40 344 42
rect 346 40 349 42
rect 341 38 349 40
rect 344 35 349 38
rect 351 46 358 48
rect 351 44 354 46
rect 356 44 358 46
rect 351 42 358 44
rect 374 46 381 51
rect 374 44 376 46
rect 378 44 381 46
rect 351 35 356 42
rect 374 41 381 44
rect 383 50 388 55
rect 396 50 401 52
rect 383 46 391 50
rect 383 44 386 46
rect 388 44 391 46
rect 383 42 391 44
rect 393 48 401 50
rect 393 46 396 48
rect 398 46 401 48
rect 393 44 401 46
rect 403 48 410 52
rect 438 49 445 55
rect 403 46 406 48
rect 408 46 410 48
rect 403 44 410 46
rect 427 46 434 49
rect 427 44 429 46
rect 431 44 434 46
rect 393 42 398 44
rect 383 41 388 42
rect 427 42 434 44
rect 429 35 434 42
rect 436 39 445 49
rect 436 37 440 39
rect 442 37 445 39
rect 436 35 445 37
rect 447 35 452 55
rect 454 48 459 55
rect 465 53 472 55
rect 465 51 467 53
rect 469 51 472 53
rect 454 46 461 48
rect 454 44 457 46
rect 459 44 461 46
rect 454 42 461 44
rect 465 46 472 51
rect 465 44 467 46
rect 469 44 472 46
rect 454 35 459 42
rect 465 41 472 44
rect 474 53 482 55
rect 474 51 477 53
rect 479 51 482 53
rect 474 41 482 51
rect 484 48 489 55
rect 539 49 546 55
rect 484 45 492 48
rect 484 43 487 45
rect 489 43 492 45
rect 484 41 492 43
rect 487 38 492 41
rect 494 42 502 48
rect 494 40 497 42
rect 499 40 502 42
rect 494 38 502 40
rect 497 35 502 38
rect 504 46 511 48
rect 504 44 507 46
rect 509 44 511 46
rect 504 42 511 44
rect 528 46 535 49
rect 528 44 530 46
rect 532 44 535 46
rect 528 42 535 44
rect 504 35 509 42
rect 530 35 535 42
rect 537 39 546 49
rect 537 37 541 39
rect 543 37 546 39
rect 537 35 546 37
rect 548 35 553 55
rect 555 48 560 55
rect 566 53 573 55
rect 566 51 568 53
rect 570 51 573 53
rect 555 46 562 48
rect 555 44 558 46
rect 560 44 562 46
rect 555 42 562 44
rect 566 46 573 51
rect 566 44 568 46
rect 570 44 573 46
rect 555 35 560 42
rect 566 41 573 44
rect 575 53 583 55
rect 575 51 578 53
rect 580 51 583 53
rect 575 41 583 51
rect 585 48 590 55
rect 638 49 645 55
rect 585 45 593 48
rect 585 43 588 45
rect 590 43 593 45
rect 585 41 593 43
rect 588 38 593 41
rect 595 42 603 48
rect 595 40 598 42
rect 600 40 603 42
rect 595 38 603 40
rect 598 35 603 38
rect 605 46 612 48
rect 605 44 608 46
rect 610 44 612 46
rect 605 42 612 44
rect 627 46 634 49
rect 627 44 629 46
rect 631 44 634 46
rect 627 42 634 44
rect 605 35 610 42
rect 629 35 634 42
rect 636 39 645 49
rect 636 37 640 39
rect 642 37 645 39
rect 636 35 645 37
rect 647 35 652 55
rect 654 48 659 55
rect 665 53 672 55
rect 665 51 667 53
rect 669 51 672 53
rect 654 46 661 48
rect 654 44 657 46
rect 659 44 661 46
rect 654 42 661 44
rect 665 46 672 51
rect 665 44 667 46
rect 669 44 672 46
rect 654 35 659 42
rect 665 41 672 44
rect 674 53 682 55
rect 674 51 677 53
rect 679 51 682 53
rect 674 41 682 51
rect 684 48 689 55
rect 684 45 692 48
rect 684 43 687 45
rect 689 43 692 45
rect 684 41 692 43
rect 687 38 692 41
rect 694 42 702 48
rect 694 40 697 42
rect 699 40 702 42
rect 694 38 702 40
rect 697 35 702 38
rect 704 46 711 48
rect 704 44 707 46
rect 709 44 711 46
rect 704 42 711 44
rect 704 35 709 42
<< pdif >>
rect 31 381 38 383
rect 31 379 33 381
rect 35 379 38 381
rect 31 374 38 379
rect 31 372 33 374
rect 35 372 38 374
rect 31 364 38 372
rect 40 375 48 383
rect 40 373 43 375
rect 45 373 48 375
rect 40 368 48 373
rect 40 366 43 368
rect 45 366 48 368
rect 40 364 48 366
rect 50 381 58 383
rect 50 379 53 381
rect 55 379 58 381
rect 50 374 58 379
rect 50 372 53 374
rect 55 372 58 374
rect 50 364 58 372
rect 52 355 58 364
rect 60 376 65 383
rect 71 381 78 383
rect 71 379 73 381
rect 75 379 78 381
rect 60 374 67 376
rect 60 372 63 374
rect 65 372 67 374
rect 60 367 67 372
rect 60 365 63 367
rect 65 365 67 367
rect 60 363 67 365
rect 71 374 78 379
rect 71 372 73 374
rect 75 372 78 374
rect 71 364 78 372
rect 80 375 88 383
rect 80 373 83 375
rect 85 373 88 375
rect 80 368 88 373
rect 80 366 83 368
rect 85 366 88 368
rect 80 364 88 366
rect 90 381 98 383
rect 90 379 93 381
rect 95 379 98 381
rect 90 374 98 379
rect 90 372 93 374
rect 95 372 98 374
rect 90 364 98 372
rect 60 355 65 363
rect 92 355 98 364
rect 100 376 105 383
rect 100 374 107 376
rect 100 372 103 374
rect 105 372 107 374
rect 100 367 107 372
rect 114 368 119 383
rect 100 365 103 367
rect 105 365 107 367
rect 100 363 107 365
rect 112 366 119 368
rect 112 364 114 366
rect 116 364 119 366
rect 100 355 105 363
rect 112 359 119 364
rect 112 357 114 359
rect 116 357 119 359
rect 112 355 119 357
rect 121 381 129 383
rect 121 379 124 381
rect 126 379 129 381
rect 121 374 129 379
rect 121 372 124 374
rect 126 372 129 374
rect 121 355 129 372
rect 131 373 139 383
rect 131 371 134 373
rect 136 371 139 373
rect 131 366 139 371
rect 131 364 134 366
rect 136 364 139 366
rect 131 355 139 364
rect 141 381 155 383
rect 141 379 146 381
rect 148 380 155 381
rect 178 381 187 383
rect 148 379 157 380
rect 141 374 157 379
rect 141 372 146 374
rect 148 372 157 374
rect 141 355 157 372
rect 159 355 164 380
rect 166 371 171 380
rect 178 379 181 381
rect 183 379 187 381
rect 178 371 187 379
rect 166 362 174 371
rect 166 360 169 362
rect 171 360 174 362
rect 166 358 174 360
rect 176 358 187 371
rect 189 371 194 383
rect 210 371 215 383
rect 189 369 196 371
rect 189 367 192 369
rect 194 367 196 369
rect 189 362 196 367
rect 189 360 192 362
rect 194 360 196 362
rect 189 358 196 360
rect 208 369 215 371
rect 208 367 210 369
rect 212 367 215 369
rect 208 362 215 367
rect 208 360 210 362
rect 212 360 215 362
rect 208 358 215 360
rect 217 381 226 383
rect 217 379 221 381
rect 223 379 226 381
rect 249 381 263 383
rect 249 380 256 381
rect 217 371 226 379
rect 233 371 238 380
rect 217 358 228 371
rect 230 362 238 371
rect 230 360 233 362
rect 235 360 238 362
rect 230 358 238 360
rect 166 355 171 358
rect 233 355 238 358
rect 240 355 245 380
rect 247 379 256 380
rect 258 379 263 381
rect 247 374 263 379
rect 247 372 256 374
rect 258 372 263 374
rect 247 355 263 372
rect 265 373 273 383
rect 265 371 268 373
rect 270 371 273 373
rect 265 366 273 371
rect 265 364 268 366
rect 270 364 273 366
rect 265 355 273 364
rect 275 381 283 383
rect 275 379 278 381
rect 280 379 283 381
rect 275 374 283 379
rect 275 372 278 374
rect 280 372 283 374
rect 275 355 283 372
rect 285 368 290 383
rect 299 376 304 383
rect 297 374 304 376
rect 297 372 299 374
rect 301 372 304 374
rect 285 366 292 368
rect 285 364 288 366
rect 290 364 292 366
rect 285 359 292 364
rect 297 367 304 372
rect 297 365 299 367
rect 301 365 304 367
rect 297 363 304 365
rect 285 357 288 359
rect 290 357 292 359
rect 285 355 292 357
rect 299 355 304 363
rect 306 381 314 383
rect 306 379 309 381
rect 311 379 314 381
rect 306 374 314 379
rect 306 372 309 374
rect 311 372 314 374
rect 306 364 314 372
rect 316 375 324 383
rect 316 373 319 375
rect 321 373 324 375
rect 316 368 324 373
rect 316 366 319 368
rect 321 366 324 368
rect 316 364 324 366
rect 326 381 333 383
rect 326 379 329 381
rect 331 379 333 381
rect 326 374 333 379
rect 339 376 344 383
rect 326 372 329 374
rect 331 372 333 374
rect 326 364 333 372
rect 337 374 344 376
rect 337 372 339 374
rect 341 372 344 374
rect 337 367 344 372
rect 337 365 339 367
rect 341 365 344 367
rect 306 355 312 364
rect 337 363 344 365
rect 339 355 344 363
rect 346 381 354 383
rect 346 379 349 381
rect 351 379 354 381
rect 346 374 354 379
rect 346 372 349 374
rect 351 372 354 374
rect 346 364 354 372
rect 356 375 364 383
rect 356 373 359 375
rect 361 373 364 375
rect 356 368 364 373
rect 356 366 359 368
rect 361 366 364 368
rect 356 364 364 366
rect 366 381 373 383
rect 366 379 369 381
rect 371 379 373 381
rect 366 374 373 379
rect 366 372 369 374
rect 371 372 373 374
rect 366 364 373 372
rect 380 371 385 383
rect 378 369 385 371
rect 378 367 380 369
rect 382 367 385 369
rect 346 355 352 364
rect 378 362 385 367
rect 378 360 380 362
rect 382 360 385 362
rect 378 358 385 360
rect 387 381 396 383
rect 387 379 391 381
rect 393 379 396 381
rect 419 381 433 383
rect 419 380 426 381
rect 387 371 396 379
rect 403 371 408 380
rect 387 358 398 371
rect 400 362 408 371
rect 400 360 403 362
rect 405 360 408 362
rect 400 358 408 360
rect 403 355 408 358
rect 410 355 415 380
rect 417 379 426 380
rect 428 379 433 381
rect 417 374 433 379
rect 417 372 426 374
rect 428 372 433 374
rect 417 355 433 372
rect 435 373 443 383
rect 435 371 438 373
rect 440 371 443 373
rect 435 366 443 371
rect 435 364 438 366
rect 440 364 443 366
rect 435 355 443 364
rect 445 381 453 383
rect 445 379 448 381
rect 450 379 453 381
rect 445 374 453 379
rect 445 372 448 374
rect 450 372 453 374
rect 445 355 453 372
rect 455 368 460 383
rect 469 376 474 383
rect 467 374 474 376
rect 467 372 469 374
rect 471 372 474 374
rect 455 366 462 368
rect 455 364 458 366
rect 460 364 462 366
rect 455 359 462 364
rect 467 367 474 372
rect 467 365 469 367
rect 471 365 474 367
rect 467 363 474 365
rect 455 357 458 359
rect 460 357 462 359
rect 455 355 462 357
rect 469 355 474 363
rect 476 381 484 383
rect 476 379 479 381
rect 481 379 484 381
rect 476 374 484 379
rect 476 372 479 374
rect 481 372 484 374
rect 476 364 484 372
rect 486 375 494 383
rect 486 373 489 375
rect 491 373 494 375
rect 486 368 494 373
rect 486 366 489 368
rect 491 366 494 368
rect 486 364 494 366
rect 496 381 503 383
rect 496 379 499 381
rect 501 379 503 381
rect 496 374 503 379
rect 509 376 514 383
rect 496 372 499 374
rect 501 372 503 374
rect 496 364 503 372
rect 507 374 514 376
rect 507 372 509 374
rect 511 372 514 374
rect 507 367 514 372
rect 507 365 509 367
rect 511 365 514 367
rect 476 355 482 364
rect 507 363 514 365
rect 509 355 514 363
rect 516 381 524 383
rect 516 379 519 381
rect 521 379 524 381
rect 516 374 524 379
rect 516 372 519 374
rect 521 372 524 374
rect 516 364 524 372
rect 526 375 534 383
rect 526 373 529 375
rect 531 373 534 375
rect 526 368 534 373
rect 526 366 529 368
rect 531 366 534 368
rect 526 364 534 366
rect 536 381 543 383
rect 536 379 539 381
rect 541 379 543 381
rect 536 374 543 379
rect 536 372 539 374
rect 541 372 543 374
rect 536 364 543 372
rect 547 381 554 383
rect 547 379 549 381
rect 551 379 554 381
rect 547 374 554 379
rect 547 372 549 374
rect 551 372 554 374
rect 547 364 554 372
rect 556 375 564 383
rect 556 373 559 375
rect 561 373 564 375
rect 556 368 564 373
rect 556 366 559 368
rect 561 366 564 368
rect 556 364 564 366
rect 566 381 574 383
rect 566 379 569 381
rect 571 379 574 381
rect 566 374 574 379
rect 566 372 569 374
rect 571 372 574 374
rect 566 364 574 372
rect 516 355 522 364
rect 568 355 574 364
rect 576 376 581 383
rect 587 381 594 383
rect 587 379 589 381
rect 591 379 594 381
rect 576 374 583 376
rect 576 372 579 374
rect 581 372 583 374
rect 576 367 583 372
rect 576 365 579 367
rect 581 365 583 367
rect 576 363 583 365
rect 587 374 594 379
rect 587 372 589 374
rect 591 372 594 374
rect 587 364 594 372
rect 596 375 604 383
rect 596 373 599 375
rect 601 373 604 375
rect 596 368 604 373
rect 596 366 599 368
rect 601 366 604 368
rect 596 364 604 366
rect 606 381 614 383
rect 606 379 609 381
rect 611 379 614 381
rect 606 374 614 379
rect 606 372 609 374
rect 611 372 614 374
rect 606 364 614 372
rect 576 355 581 363
rect 608 355 614 364
rect 616 376 621 383
rect 616 374 623 376
rect 616 372 619 374
rect 621 372 623 374
rect 616 367 623 372
rect 630 368 635 383
rect 616 365 619 367
rect 621 365 623 367
rect 616 363 623 365
rect 628 366 635 368
rect 628 364 630 366
rect 632 364 635 366
rect 616 355 621 363
rect 628 359 635 364
rect 628 357 630 359
rect 632 357 635 359
rect 628 355 635 357
rect 637 381 645 383
rect 637 379 640 381
rect 642 379 645 381
rect 637 374 645 379
rect 637 372 640 374
rect 642 372 645 374
rect 637 355 645 372
rect 647 373 655 383
rect 647 371 650 373
rect 652 371 655 373
rect 647 366 655 371
rect 647 364 650 366
rect 652 364 655 366
rect 647 355 655 364
rect 657 381 671 383
rect 657 379 662 381
rect 664 380 671 381
rect 694 381 703 383
rect 664 379 673 380
rect 657 374 673 379
rect 657 372 662 374
rect 664 372 673 374
rect 657 355 673 372
rect 675 355 680 380
rect 682 371 687 380
rect 694 379 697 381
rect 699 379 703 381
rect 694 371 703 379
rect 682 362 690 371
rect 682 360 685 362
rect 687 360 690 362
rect 682 358 690 360
rect 692 358 703 371
rect 705 371 710 383
rect 705 369 712 371
rect 705 367 708 369
rect 710 367 712 369
rect 705 362 712 367
rect 705 360 708 362
rect 710 360 712 362
rect 705 358 712 360
rect 682 355 687 358
rect 52 270 58 279
rect 31 262 38 270
rect 31 260 33 262
rect 35 260 38 262
rect 31 255 38 260
rect 31 253 33 255
rect 35 253 38 255
rect 31 251 38 253
rect 40 268 48 270
rect 40 266 43 268
rect 45 266 48 268
rect 40 261 48 266
rect 40 259 43 261
rect 45 259 48 261
rect 40 251 48 259
rect 50 262 58 270
rect 50 260 53 262
rect 55 260 58 262
rect 50 255 58 260
rect 50 253 53 255
rect 55 253 58 255
rect 50 251 58 253
rect 60 271 65 279
rect 60 269 67 271
rect 92 270 98 279
rect 60 267 63 269
rect 65 267 67 269
rect 60 262 67 267
rect 60 260 63 262
rect 65 260 67 262
rect 60 258 67 260
rect 71 262 78 270
rect 71 260 73 262
rect 75 260 78 262
rect 60 251 65 258
rect 71 255 78 260
rect 71 253 73 255
rect 75 253 78 255
rect 71 251 78 253
rect 80 268 88 270
rect 80 266 83 268
rect 85 266 88 268
rect 80 261 88 266
rect 80 259 83 261
rect 85 259 88 261
rect 80 251 88 259
rect 90 262 98 270
rect 90 260 93 262
rect 95 260 98 262
rect 90 255 98 260
rect 90 253 93 255
rect 95 253 98 255
rect 90 251 98 253
rect 100 271 105 279
rect 112 277 119 279
rect 112 275 114 277
rect 116 275 119 277
rect 100 269 107 271
rect 100 267 103 269
rect 105 267 107 269
rect 100 262 107 267
rect 112 266 119 275
rect 100 260 103 262
rect 105 260 107 262
rect 100 258 107 260
rect 100 251 105 258
rect 114 251 119 266
rect 121 262 129 279
rect 121 260 124 262
rect 126 260 129 262
rect 121 255 129 260
rect 121 253 124 255
rect 126 253 129 255
rect 121 251 129 253
rect 131 270 139 279
rect 131 268 134 270
rect 136 268 139 270
rect 131 263 139 268
rect 131 261 134 263
rect 136 261 139 263
rect 131 251 139 261
rect 141 262 157 279
rect 141 260 146 262
rect 148 260 157 262
rect 141 255 157 260
rect 141 253 146 255
rect 148 254 157 255
rect 159 254 164 279
rect 166 276 171 279
rect 233 276 238 279
rect 166 274 174 276
rect 166 272 169 274
rect 171 272 174 274
rect 166 263 174 272
rect 176 263 187 276
rect 166 254 171 263
rect 178 255 187 263
rect 148 253 155 254
rect 141 251 155 253
rect 178 253 181 255
rect 183 253 187 255
rect 178 251 187 253
rect 189 274 196 276
rect 189 272 192 274
rect 194 272 196 274
rect 189 267 196 272
rect 189 265 192 267
rect 194 265 196 267
rect 189 263 196 265
rect 208 274 215 276
rect 208 272 210 274
rect 212 272 215 274
rect 208 267 215 272
rect 208 265 210 267
rect 212 265 215 267
rect 208 263 215 265
rect 189 251 194 263
rect 210 251 215 263
rect 217 263 228 276
rect 230 274 238 276
rect 230 272 233 274
rect 235 272 238 274
rect 230 263 238 272
rect 217 255 226 263
rect 217 253 221 255
rect 223 253 226 255
rect 233 254 238 263
rect 240 254 245 279
rect 247 262 263 279
rect 247 260 256 262
rect 258 260 263 262
rect 247 255 263 260
rect 247 254 256 255
rect 217 251 226 253
rect 249 253 256 254
rect 258 253 263 255
rect 249 251 263 253
rect 265 270 273 279
rect 265 268 268 270
rect 270 268 273 270
rect 265 263 273 268
rect 265 261 268 263
rect 270 261 273 263
rect 265 251 273 261
rect 275 262 283 279
rect 275 260 278 262
rect 280 260 283 262
rect 275 255 283 260
rect 275 253 278 255
rect 280 253 283 255
rect 275 251 283 253
rect 285 277 292 279
rect 285 275 288 277
rect 290 275 292 277
rect 285 270 292 275
rect 299 271 304 279
rect 285 268 288 270
rect 290 268 292 270
rect 285 266 292 268
rect 297 269 304 271
rect 297 267 299 269
rect 301 267 304 269
rect 285 251 290 266
rect 297 262 304 267
rect 297 260 299 262
rect 301 260 304 262
rect 297 258 304 260
rect 299 251 304 258
rect 306 270 312 279
rect 339 271 344 279
rect 306 262 314 270
rect 306 260 309 262
rect 311 260 314 262
rect 306 255 314 260
rect 306 253 309 255
rect 311 253 314 255
rect 306 251 314 253
rect 316 268 324 270
rect 316 266 319 268
rect 321 266 324 268
rect 316 261 324 266
rect 316 259 319 261
rect 321 259 324 261
rect 316 251 324 259
rect 326 262 333 270
rect 326 260 329 262
rect 331 260 333 262
rect 326 255 333 260
rect 337 269 344 271
rect 337 267 339 269
rect 341 267 344 269
rect 337 262 344 267
rect 337 260 339 262
rect 341 260 344 262
rect 337 258 344 260
rect 326 253 329 255
rect 331 253 333 255
rect 326 251 333 253
rect 339 251 344 258
rect 346 270 352 279
rect 403 276 408 279
rect 378 274 385 276
rect 378 272 380 274
rect 382 272 385 274
rect 346 262 354 270
rect 346 260 349 262
rect 351 260 354 262
rect 346 255 354 260
rect 346 253 349 255
rect 351 253 354 255
rect 346 251 354 253
rect 356 268 364 270
rect 356 266 359 268
rect 361 266 364 268
rect 356 261 364 266
rect 356 259 359 261
rect 361 259 364 261
rect 356 251 364 259
rect 366 262 373 270
rect 378 267 385 272
rect 378 265 380 267
rect 382 265 385 267
rect 378 263 385 265
rect 366 260 369 262
rect 371 260 373 262
rect 366 255 373 260
rect 366 253 369 255
rect 371 253 373 255
rect 366 251 373 253
rect 380 251 385 263
rect 387 263 398 276
rect 400 274 408 276
rect 400 272 403 274
rect 405 272 408 274
rect 400 263 408 272
rect 387 255 396 263
rect 387 253 391 255
rect 393 253 396 255
rect 403 254 408 263
rect 410 254 415 279
rect 417 262 433 279
rect 417 260 426 262
rect 428 260 433 262
rect 417 255 433 260
rect 417 254 426 255
rect 387 251 396 253
rect 419 253 426 254
rect 428 253 433 255
rect 419 251 433 253
rect 435 270 443 279
rect 435 268 438 270
rect 440 268 443 270
rect 435 263 443 268
rect 435 261 438 263
rect 440 261 443 263
rect 435 251 443 261
rect 445 262 453 279
rect 445 260 448 262
rect 450 260 453 262
rect 445 255 453 260
rect 445 253 448 255
rect 450 253 453 255
rect 445 251 453 253
rect 455 277 462 279
rect 455 275 458 277
rect 460 275 462 277
rect 455 270 462 275
rect 469 271 474 279
rect 455 268 458 270
rect 460 268 462 270
rect 455 266 462 268
rect 467 269 474 271
rect 467 267 469 269
rect 471 267 474 269
rect 455 251 460 266
rect 467 262 474 267
rect 467 260 469 262
rect 471 260 474 262
rect 467 258 474 260
rect 469 251 474 258
rect 476 270 482 279
rect 509 271 514 279
rect 476 262 484 270
rect 476 260 479 262
rect 481 260 484 262
rect 476 255 484 260
rect 476 253 479 255
rect 481 253 484 255
rect 476 251 484 253
rect 486 268 494 270
rect 486 266 489 268
rect 491 266 494 268
rect 486 261 494 266
rect 486 259 489 261
rect 491 259 494 261
rect 486 251 494 259
rect 496 262 503 270
rect 496 260 499 262
rect 501 260 503 262
rect 496 255 503 260
rect 507 269 514 271
rect 507 267 509 269
rect 511 267 514 269
rect 507 262 514 267
rect 507 260 509 262
rect 511 260 514 262
rect 507 258 514 260
rect 496 253 499 255
rect 501 253 503 255
rect 496 251 503 253
rect 509 251 514 258
rect 516 270 522 279
rect 568 270 574 279
rect 516 262 524 270
rect 516 260 519 262
rect 521 260 524 262
rect 516 255 524 260
rect 516 253 519 255
rect 521 253 524 255
rect 516 251 524 253
rect 526 268 534 270
rect 526 266 529 268
rect 531 266 534 268
rect 526 261 534 266
rect 526 259 529 261
rect 531 259 534 261
rect 526 251 534 259
rect 536 262 543 270
rect 536 260 539 262
rect 541 260 543 262
rect 536 255 543 260
rect 536 253 539 255
rect 541 253 543 255
rect 536 251 543 253
rect 547 262 554 270
rect 547 260 549 262
rect 551 260 554 262
rect 547 255 554 260
rect 547 253 549 255
rect 551 253 554 255
rect 547 251 554 253
rect 556 268 564 270
rect 556 266 559 268
rect 561 266 564 268
rect 556 261 564 266
rect 556 259 559 261
rect 561 259 564 261
rect 556 251 564 259
rect 566 262 574 270
rect 566 260 569 262
rect 571 260 574 262
rect 566 255 574 260
rect 566 253 569 255
rect 571 253 574 255
rect 566 251 574 253
rect 576 271 581 279
rect 576 269 583 271
rect 608 270 614 279
rect 576 267 579 269
rect 581 267 583 269
rect 576 262 583 267
rect 576 260 579 262
rect 581 260 583 262
rect 576 258 583 260
rect 587 262 594 270
rect 587 260 589 262
rect 591 260 594 262
rect 576 251 581 258
rect 587 255 594 260
rect 587 253 589 255
rect 591 253 594 255
rect 587 251 594 253
rect 596 268 604 270
rect 596 266 599 268
rect 601 266 604 268
rect 596 261 604 266
rect 596 259 599 261
rect 601 259 604 261
rect 596 251 604 259
rect 606 262 614 270
rect 606 260 609 262
rect 611 260 614 262
rect 606 255 614 260
rect 606 253 609 255
rect 611 253 614 255
rect 606 251 614 253
rect 616 271 621 279
rect 628 277 635 279
rect 628 275 630 277
rect 632 275 635 277
rect 616 269 623 271
rect 616 267 619 269
rect 621 267 623 269
rect 616 262 623 267
rect 628 270 635 275
rect 628 268 630 270
rect 632 268 635 270
rect 628 266 635 268
rect 616 260 619 262
rect 621 260 623 262
rect 616 258 623 260
rect 616 251 621 258
rect 630 251 635 266
rect 637 262 645 279
rect 637 260 640 262
rect 642 260 645 262
rect 637 255 645 260
rect 637 253 640 255
rect 642 253 645 255
rect 637 251 645 253
rect 647 270 655 279
rect 647 268 650 270
rect 652 268 655 270
rect 647 263 655 268
rect 647 261 650 263
rect 652 261 655 263
rect 647 251 655 261
rect 657 262 673 279
rect 657 260 662 262
rect 664 260 673 262
rect 657 255 673 260
rect 657 253 662 255
rect 664 254 673 255
rect 675 254 680 279
rect 682 276 687 279
rect 682 274 690 276
rect 682 272 685 274
rect 687 272 690 274
rect 682 263 690 272
rect 692 263 703 276
rect 682 254 687 263
rect 694 255 703 263
rect 664 253 671 254
rect 657 251 671 253
rect 694 253 697 255
rect 699 253 703 255
rect 694 251 703 253
rect 705 274 712 276
rect 705 272 708 274
rect 710 272 712 274
rect 705 267 712 272
rect 705 265 708 267
rect 710 265 712 267
rect 705 263 712 265
rect 705 251 710 263
rect 42 240 49 242
rect 42 239 44 240
rect 33 233 38 239
rect 31 231 38 233
rect 31 229 33 231
rect 35 229 38 231
rect 31 224 38 229
rect 31 222 33 224
rect 35 222 38 224
rect 31 220 38 222
rect 33 211 38 220
rect 40 238 44 239
rect 46 239 49 240
rect 46 238 51 239
rect 40 211 51 238
rect 53 211 58 239
rect 60 233 65 239
rect 60 231 67 233
rect 60 229 63 231
rect 65 229 67 231
rect 60 227 67 229
rect 60 211 65 227
rect 74 224 79 239
rect 72 222 79 224
rect 72 220 74 222
rect 76 220 79 222
rect 72 215 79 220
rect 72 213 74 215
rect 76 213 79 215
rect 72 211 79 213
rect 81 237 89 239
rect 81 235 84 237
rect 86 235 89 237
rect 81 230 89 235
rect 81 228 84 230
rect 86 228 89 230
rect 81 211 89 228
rect 91 229 99 239
rect 91 227 94 229
rect 96 227 99 229
rect 91 222 99 227
rect 91 220 94 222
rect 96 220 99 222
rect 91 211 99 220
rect 101 237 115 239
rect 101 235 106 237
rect 108 236 115 237
rect 138 237 147 239
rect 108 235 117 236
rect 101 230 117 235
rect 101 228 106 230
rect 108 228 117 230
rect 101 211 117 228
rect 119 211 124 236
rect 126 227 131 236
rect 138 235 141 237
rect 143 235 147 237
rect 138 227 147 235
rect 126 218 134 227
rect 126 216 129 218
rect 131 216 134 218
rect 126 214 134 216
rect 136 214 147 227
rect 149 227 154 239
rect 149 225 156 227
rect 149 223 152 225
rect 154 223 156 225
rect 175 224 180 239
rect 149 218 156 223
rect 149 216 152 218
rect 154 216 156 218
rect 149 214 156 216
rect 173 222 180 224
rect 173 220 175 222
rect 177 220 180 222
rect 173 215 180 220
rect 126 211 131 214
rect 173 213 175 215
rect 177 213 180 215
rect 173 211 180 213
rect 182 237 190 239
rect 182 235 185 237
rect 187 235 190 237
rect 182 230 190 235
rect 182 228 185 230
rect 187 228 190 230
rect 182 211 190 228
rect 192 229 200 239
rect 192 227 195 229
rect 197 227 200 229
rect 192 222 200 227
rect 192 220 195 222
rect 197 220 200 222
rect 192 211 200 220
rect 202 237 216 239
rect 202 235 207 237
rect 209 236 216 237
rect 239 237 248 239
rect 209 235 218 236
rect 202 230 218 235
rect 202 228 207 230
rect 209 228 218 230
rect 202 211 218 228
rect 220 211 225 236
rect 227 227 232 236
rect 239 235 242 237
rect 244 235 248 237
rect 239 227 248 235
rect 227 218 235 227
rect 227 216 230 218
rect 232 216 235 218
rect 227 214 235 216
rect 237 214 248 227
rect 250 227 255 239
rect 250 225 257 227
rect 250 223 253 225
rect 255 223 257 225
rect 277 224 282 239
rect 250 218 257 223
rect 250 216 253 218
rect 255 216 257 218
rect 250 214 257 216
rect 275 222 282 224
rect 275 220 277 222
rect 279 220 282 222
rect 275 215 282 220
rect 227 211 232 214
rect 275 213 277 215
rect 279 213 282 215
rect 275 211 282 213
rect 284 237 292 239
rect 284 235 287 237
rect 289 235 292 237
rect 284 230 292 235
rect 284 228 287 230
rect 289 228 292 230
rect 284 211 292 228
rect 294 229 302 239
rect 294 227 297 229
rect 299 227 302 229
rect 294 222 302 227
rect 294 220 297 222
rect 299 220 302 222
rect 294 211 302 220
rect 304 237 318 239
rect 304 235 309 237
rect 311 236 318 237
rect 386 240 393 242
rect 386 239 388 240
rect 341 237 350 239
rect 311 235 320 236
rect 304 230 320 235
rect 304 228 309 230
rect 311 228 320 230
rect 304 211 320 228
rect 322 211 327 236
rect 329 227 334 236
rect 341 235 344 237
rect 346 235 350 237
rect 341 227 350 235
rect 329 218 337 227
rect 329 216 332 218
rect 334 216 337 218
rect 329 214 337 216
rect 339 214 350 227
rect 352 227 357 239
rect 377 233 382 239
rect 375 231 382 233
rect 375 229 377 231
rect 379 229 382 231
rect 352 225 359 227
rect 352 223 355 225
rect 357 223 359 225
rect 352 218 359 223
rect 375 224 382 229
rect 375 222 377 224
rect 379 222 382 224
rect 375 220 382 222
rect 352 216 355 218
rect 357 216 359 218
rect 352 214 359 216
rect 329 211 334 214
rect 377 211 382 220
rect 384 238 388 239
rect 390 239 393 240
rect 390 238 395 239
rect 384 211 395 238
rect 397 211 402 239
rect 404 233 409 239
rect 404 231 411 233
rect 404 229 407 231
rect 409 229 411 231
rect 404 227 411 229
rect 404 211 409 227
rect 430 224 435 239
rect 428 222 435 224
rect 428 220 430 222
rect 432 220 435 222
rect 428 215 435 220
rect 428 213 430 215
rect 432 213 435 215
rect 428 211 435 213
rect 437 237 445 239
rect 437 235 440 237
rect 442 235 445 237
rect 437 230 445 235
rect 437 228 440 230
rect 442 228 445 230
rect 437 211 445 228
rect 447 229 455 239
rect 447 227 450 229
rect 452 227 455 229
rect 447 222 455 227
rect 447 220 450 222
rect 452 220 455 222
rect 447 211 455 220
rect 457 237 471 239
rect 457 235 462 237
rect 464 236 471 237
rect 494 237 503 239
rect 464 235 473 236
rect 457 230 473 235
rect 457 228 462 230
rect 464 228 473 230
rect 457 211 473 228
rect 475 211 480 236
rect 482 227 487 236
rect 494 235 497 237
rect 499 235 503 237
rect 494 227 503 235
rect 482 218 490 227
rect 482 216 485 218
rect 487 216 490 218
rect 482 214 490 216
rect 492 214 503 227
rect 505 227 510 239
rect 505 225 512 227
rect 505 223 508 225
rect 510 223 512 225
rect 531 224 536 239
rect 505 218 512 223
rect 505 216 508 218
rect 510 216 512 218
rect 505 214 512 216
rect 529 222 536 224
rect 529 220 531 222
rect 533 220 536 222
rect 529 215 536 220
rect 482 211 487 214
rect 529 213 531 215
rect 533 213 536 215
rect 529 211 536 213
rect 538 237 546 239
rect 538 235 541 237
rect 543 235 546 237
rect 538 230 546 235
rect 538 228 541 230
rect 543 228 546 230
rect 538 211 546 228
rect 548 229 556 239
rect 548 227 551 229
rect 553 227 556 229
rect 548 222 556 227
rect 548 220 551 222
rect 553 220 556 222
rect 548 211 556 220
rect 558 237 572 239
rect 558 235 563 237
rect 565 236 572 237
rect 595 237 604 239
rect 565 235 574 236
rect 558 230 574 235
rect 558 228 563 230
rect 565 228 574 230
rect 558 211 574 228
rect 576 211 581 236
rect 583 227 588 236
rect 595 235 598 237
rect 600 235 604 237
rect 595 227 604 235
rect 583 218 591 227
rect 583 216 586 218
rect 588 216 591 218
rect 583 214 591 216
rect 593 214 604 227
rect 606 227 611 239
rect 606 225 613 227
rect 606 223 609 225
rect 611 223 613 225
rect 630 224 635 239
rect 606 218 613 223
rect 606 216 609 218
rect 611 216 613 218
rect 606 214 613 216
rect 628 222 635 224
rect 628 220 630 222
rect 632 220 635 222
rect 628 215 635 220
rect 583 211 588 214
rect 628 213 630 215
rect 632 213 635 215
rect 628 211 635 213
rect 637 237 645 239
rect 637 235 640 237
rect 642 235 645 237
rect 637 230 645 235
rect 637 228 640 230
rect 642 228 645 230
rect 637 211 645 228
rect 647 229 655 239
rect 647 227 650 229
rect 652 227 655 229
rect 647 222 655 227
rect 647 220 650 222
rect 652 220 655 222
rect 647 211 655 220
rect 657 237 671 239
rect 657 235 662 237
rect 664 236 671 237
rect 694 237 703 239
rect 664 235 673 236
rect 657 230 673 235
rect 657 228 662 230
rect 664 228 673 230
rect 657 211 673 228
rect 675 211 680 236
rect 682 227 687 236
rect 694 235 697 237
rect 699 235 703 237
rect 694 227 703 235
rect 682 218 690 227
rect 682 216 685 218
rect 687 216 690 218
rect 682 214 690 216
rect 692 214 703 227
rect 705 227 710 239
rect 705 225 712 227
rect 705 223 708 225
rect 710 223 712 225
rect 705 218 712 223
rect 705 216 708 218
rect 710 216 712 218
rect 705 214 712 216
rect 682 211 687 214
rect 33 133 40 135
rect 33 131 35 133
rect 37 131 40 133
rect 33 126 40 131
rect 33 124 35 126
rect 37 124 40 126
rect 33 122 40 124
rect 35 107 40 122
rect 42 118 50 135
rect 42 116 45 118
rect 47 116 50 118
rect 42 111 50 116
rect 42 109 45 111
rect 47 109 50 111
rect 42 107 50 109
rect 52 126 60 135
rect 52 124 55 126
rect 57 124 60 126
rect 52 119 60 124
rect 52 117 55 119
rect 57 117 60 119
rect 52 107 60 117
rect 62 118 78 135
rect 62 116 67 118
rect 69 116 78 118
rect 62 111 78 116
rect 62 109 67 111
rect 69 110 78 111
rect 80 110 85 135
rect 87 132 92 135
rect 87 130 95 132
rect 87 128 90 130
rect 92 128 95 130
rect 87 119 95 128
rect 97 119 108 132
rect 87 110 92 119
rect 99 111 108 119
rect 69 109 76 110
rect 62 107 76 109
rect 99 109 102 111
rect 104 109 108 111
rect 99 107 108 109
rect 110 130 117 132
rect 110 128 113 130
rect 115 128 117 130
rect 110 123 117 128
rect 123 126 128 135
rect 110 121 113 123
rect 115 121 117 123
rect 110 119 117 121
rect 121 124 128 126
rect 121 122 123 124
rect 125 122 128 124
rect 110 107 115 119
rect 121 117 128 122
rect 121 115 123 117
rect 125 115 128 117
rect 121 113 128 115
rect 123 107 128 113
rect 130 108 141 135
rect 130 107 134 108
rect 132 106 134 107
rect 136 107 141 108
rect 143 107 148 135
rect 150 119 155 135
rect 174 133 181 135
rect 174 131 176 133
rect 178 131 181 133
rect 174 126 181 131
rect 174 124 176 126
rect 178 124 181 126
rect 174 122 181 124
rect 150 117 157 119
rect 150 115 153 117
rect 155 115 157 117
rect 150 113 157 115
rect 150 107 155 113
rect 176 107 181 122
rect 183 118 191 135
rect 183 116 186 118
rect 188 116 191 118
rect 183 111 191 116
rect 183 109 186 111
rect 188 109 191 111
rect 183 107 191 109
rect 193 126 201 135
rect 193 124 196 126
rect 198 124 201 126
rect 193 119 201 124
rect 193 117 196 119
rect 198 117 201 119
rect 193 107 201 117
rect 203 118 219 135
rect 203 116 208 118
rect 210 116 219 118
rect 203 111 219 116
rect 203 109 208 111
rect 210 110 219 111
rect 221 110 226 135
rect 228 132 233 135
rect 299 132 304 135
rect 228 130 236 132
rect 228 128 231 130
rect 233 128 236 130
rect 228 119 236 128
rect 238 119 249 132
rect 228 110 233 119
rect 240 111 249 119
rect 210 109 217 110
rect 203 107 217 109
rect 136 106 139 107
rect 132 104 139 106
rect 240 109 243 111
rect 245 109 249 111
rect 240 107 249 109
rect 251 130 258 132
rect 251 128 254 130
rect 256 128 258 130
rect 251 123 258 128
rect 251 121 254 123
rect 256 121 258 123
rect 251 119 258 121
rect 274 130 281 132
rect 274 128 276 130
rect 278 128 281 130
rect 274 123 281 128
rect 274 121 276 123
rect 278 121 281 123
rect 274 119 281 121
rect 251 107 256 119
rect 276 107 281 119
rect 283 119 294 132
rect 296 130 304 132
rect 296 128 299 130
rect 301 128 304 130
rect 296 119 304 128
rect 283 111 292 119
rect 283 109 287 111
rect 289 109 292 111
rect 299 110 304 119
rect 306 110 311 135
rect 313 118 329 135
rect 313 116 322 118
rect 324 116 329 118
rect 313 111 329 116
rect 313 110 322 111
rect 283 107 292 109
rect 315 109 322 110
rect 324 109 329 111
rect 315 107 329 109
rect 331 126 339 135
rect 331 124 334 126
rect 336 124 339 126
rect 331 119 339 124
rect 331 117 334 119
rect 336 117 339 119
rect 331 107 339 117
rect 341 118 349 135
rect 341 116 344 118
rect 346 116 349 118
rect 341 111 349 116
rect 341 109 344 111
rect 346 109 349 111
rect 341 107 349 109
rect 351 133 358 135
rect 351 131 354 133
rect 356 131 358 133
rect 351 126 358 131
rect 377 126 382 135
rect 351 124 354 126
rect 356 124 358 126
rect 351 122 358 124
rect 375 124 382 126
rect 375 122 377 124
rect 379 122 382 124
rect 351 107 356 122
rect 375 117 382 122
rect 375 115 377 117
rect 379 115 382 117
rect 375 113 382 115
rect 377 107 382 113
rect 384 108 395 135
rect 384 107 388 108
rect 386 106 388 107
rect 390 107 395 108
rect 397 107 402 135
rect 404 119 409 135
rect 428 133 435 135
rect 428 131 430 133
rect 432 131 435 133
rect 428 126 435 131
rect 428 124 430 126
rect 432 124 435 126
rect 428 122 435 124
rect 404 117 411 119
rect 404 115 407 117
rect 409 115 411 117
rect 404 113 411 115
rect 404 107 409 113
rect 430 107 435 122
rect 437 118 445 135
rect 437 116 440 118
rect 442 116 445 118
rect 437 111 445 116
rect 437 109 440 111
rect 442 109 445 111
rect 437 107 445 109
rect 447 126 455 135
rect 447 124 450 126
rect 452 124 455 126
rect 447 119 455 124
rect 447 117 450 119
rect 452 117 455 119
rect 447 107 455 117
rect 457 118 473 135
rect 457 116 462 118
rect 464 116 473 118
rect 457 111 473 116
rect 457 109 462 111
rect 464 110 473 111
rect 475 110 480 135
rect 482 132 487 135
rect 529 133 536 135
rect 482 130 490 132
rect 482 128 485 130
rect 487 128 490 130
rect 482 119 490 128
rect 492 119 503 132
rect 482 110 487 119
rect 494 111 503 119
rect 464 109 471 110
rect 457 107 471 109
rect 390 106 393 107
rect 386 104 393 106
rect 494 109 497 111
rect 499 109 503 111
rect 494 107 503 109
rect 505 130 512 132
rect 505 128 508 130
rect 510 128 512 130
rect 505 123 512 128
rect 505 121 508 123
rect 510 121 512 123
rect 529 131 531 133
rect 533 131 536 133
rect 529 126 536 131
rect 529 124 531 126
rect 533 124 536 126
rect 529 122 536 124
rect 505 119 512 121
rect 505 107 510 119
rect 531 107 536 122
rect 538 118 546 135
rect 538 116 541 118
rect 543 116 546 118
rect 538 111 546 116
rect 538 109 541 111
rect 543 109 546 111
rect 538 107 546 109
rect 548 126 556 135
rect 548 124 551 126
rect 553 124 556 126
rect 548 119 556 124
rect 548 117 551 119
rect 553 117 556 119
rect 548 107 556 117
rect 558 118 574 135
rect 558 116 563 118
rect 565 116 574 118
rect 558 111 574 116
rect 558 109 563 111
rect 565 110 574 111
rect 576 110 581 135
rect 583 132 588 135
rect 628 133 635 135
rect 583 130 591 132
rect 583 128 586 130
rect 588 128 591 130
rect 583 119 591 128
rect 593 119 604 132
rect 583 110 588 119
rect 595 111 604 119
rect 565 109 572 110
rect 558 107 572 109
rect 595 109 598 111
rect 600 109 604 111
rect 595 107 604 109
rect 606 130 613 132
rect 606 128 609 130
rect 611 128 613 130
rect 606 123 613 128
rect 606 121 609 123
rect 611 121 613 123
rect 628 131 630 133
rect 632 131 635 133
rect 628 126 635 131
rect 628 124 630 126
rect 632 124 635 126
rect 628 122 635 124
rect 606 119 613 121
rect 606 107 611 119
rect 630 107 635 122
rect 637 118 645 135
rect 637 116 640 118
rect 642 116 645 118
rect 637 111 645 116
rect 637 109 640 111
rect 642 109 645 111
rect 637 107 645 109
rect 647 126 655 135
rect 647 124 650 126
rect 652 124 655 126
rect 647 119 655 124
rect 647 117 650 119
rect 652 117 655 119
rect 647 107 655 117
rect 657 118 673 135
rect 657 116 662 118
rect 664 116 673 118
rect 657 111 673 116
rect 657 109 662 111
rect 664 110 673 111
rect 675 110 680 135
rect 682 132 687 135
rect 682 130 690 132
rect 682 128 685 130
rect 687 128 690 130
rect 682 119 690 128
rect 692 119 703 132
rect 682 110 687 119
rect 694 111 703 119
rect 664 109 671 110
rect 657 107 671 109
rect 694 109 697 111
rect 699 109 703 111
rect 694 107 703 109
rect 705 130 712 132
rect 705 128 708 130
rect 710 128 712 130
rect 705 123 712 128
rect 705 121 708 123
rect 710 121 712 123
rect 705 119 712 121
rect 705 107 710 119
rect 42 96 49 98
rect 42 95 44 96
rect 33 89 38 95
rect 31 87 38 89
rect 31 85 33 87
rect 35 85 38 87
rect 31 80 38 85
rect 31 78 33 80
rect 35 78 38 80
rect 31 76 38 78
rect 33 67 38 76
rect 40 94 44 95
rect 46 95 49 96
rect 46 94 51 95
rect 40 67 51 94
rect 53 67 58 95
rect 60 89 65 95
rect 60 87 67 89
rect 60 85 63 87
rect 65 85 67 87
rect 60 83 67 85
rect 60 67 65 83
rect 74 80 79 95
rect 72 78 79 80
rect 72 76 74 78
rect 76 76 79 78
rect 72 71 79 76
rect 72 69 74 71
rect 76 69 79 71
rect 72 67 79 69
rect 81 93 89 95
rect 81 91 84 93
rect 86 91 89 93
rect 81 86 89 91
rect 81 84 84 86
rect 86 84 89 86
rect 81 67 89 84
rect 91 85 99 95
rect 91 83 94 85
rect 96 83 99 85
rect 91 78 99 83
rect 91 76 94 78
rect 96 76 99 78
rect 91 67 99 76
rect 101 93 115 95
rect 101 91 106 93
rect 108 92 115 93
rect 138 93 147 95
rect 108 91 117 92
rect 101 86 117 91
rect 101 84 106 86
rect 108 84 117 86
rect 101 67 117 84
rect 119 67 124 92
rect 126 83 131 92
rect 138 91 141 93
rect 143 91 147 93
rect 138 83 147 91
rect 126 74 134 83
rect 126 72 129 74
rect 131 72 134 74
rect 126 70 134 72
rect 136 70 147 83
rect 149 83 154 95
rect 149 81 156 83
rect 149 79 152 81
rect 154 79 156 81
rect 175 80 180 95
rect 149 74 156 79
rect 149 72 152 74
rect 154 72 156 74
rect 149 70 156 72
rect 173 78 180 80
rect 173 76 175 78
rect 177 76 180 78
rect 173 71 180 76
rect 126 67 131 70
rect 173 69 175 71
rect 177 69 180 71
rect 173 67 180 69
rect 182 93 190 95
rect 182 91 185 93
rect 187 91 190 93
rect 182 86 190 91
rect 182 84 185 86
rect 187 84 190 86
rect 182 67 190 84
rect 192 85 200 95
rect 192 83 195 85
rect 197 83 200 85
rect 192 78 200 83
rect 192 76 195 78
rect 197 76 200 78
rect 192 67 200 76
rect 202 93 216 95
rect 202 91 207 93
rect 209 92 216 93
rect 239 93 248 95
rect 209 91 218 92
rect 202 86 218 91
rect 202 84 207 86
rect 209 84 218 86
rect 202 67 218 84
rect 220 67 225 92
rect 227 83 232 92
rect 239 91 242 93
rect 244 91 248 93
rect 239 83 248 91
rect 227 74 235 83
rect 227 72 230 74
rect 232 72 235 74
rect 227 70 235 72
rect 237 70 248 83
rect 250 83 255 95
rect 250 81 257 83
rect 250 79 253 81
rect 255 79 257 81
rect 276 80 281 95
rect 250 74 257 79
rect 250 72 253 74
rect 255 72 257 74
rect 250 70 257 72
rect 274 78 281 80
rect 274 76 276 78
rect 278 76 281 78
rect 274 71 281 76
rect 227 67 232 70
rect 274 69 276 71
rect 278 69 281 71
rect 274 67 281 69
rect 283 93 291 95
rect 283 91 286 93
rect 288 91 291 93
rect 283 86 291 91
rect 283 84 286 86
rect 288 84 291 86
rect 283 67 291 84
rect 293 85 301 95
rect 293 83 296 85
rect 298 83 301 85
rect 293 78 301 83
rect 293 76 296 78
rect 298 76 301 78
rect 293 67 301 76
rect 303 93 317 95
rect 303 91 308 93
rect 310 92 317 93
rect 385 96 392 98
rect 385 95 387 96
rect 340 93 349 95
rect 310 91 319 92
rect 303 86 319 91
rect 303 84 308 86
rect 310 84 319 86
rect 303 67 319 84
rect 321 67 326 92
rect 328 83 333 92
rect 340 91 343 93
rect 345 91 349 93
rect 340 83 349 91
rect 328 74 336 83
rect 328 72 331 74
rect 333 72 336 74
rect 328 70 336 72
rect 338 70 349 83
rect 351 83 356 95
rect 376 89 381 95
rect 374 87 381 89
rect 374 85 376 87
rect 378 85 381 87
rect 351 81 358 83
rect 351 79 354 81
rect 356 79 358 81
rect 351 74 358 79
rect 374 80 381 85
rect 374 78 376 80
rect 378 78 381 80
rect 374 76 381 78
rect 351 72 354 74
rect 356 72 358 74
rect 351 70 358 72
rect 328 67 333 70
rect 376 67 381 76
rect 383 94 387 95
rect 389 95 392 96
rect 389 94 394 95
rect 383 67 394 94
rect 396 67 401 95
rect 403 89 408 95
rect 403 87 410 89
rect 403 85 406 87
rect 408 85 410 87
rect 403 83 410 85
rect 403 67 408 83
rect 429 80 434 95
rect 427 78 434 80
rect 427 76 429 78
rect 431 76 434 78
rect 427 71 434 76
rect 427 69 429 71
rect 431 69 434 71
rect 427 67 434 69
rect 436 93 444 95
rect 436 91 439 93
rect 441 91 444 93
rect 436 86 444 91
rect 436 84 439 86
rect 441 84 444 86
rect 436 67 444 84
rect 446 85 454 95
rect 446 83 449 85
rect 451 83 454 85
rect 446 78 454 83
rect 446 76 449 78
rect 451 76 454 78
rect 446 67 454 76
rect 456 93 470 95
rect 456 91 461 93
rect 463 92 470 93
rect 493 93 502 95
rect 463 91 472 92
rect 456 86 472 91
rect 456 84 461 86
rect 463 84 472 86
rect 456 67 472 84
rect 474 67 479 92
rect 481 83 486 92
rect 493 91 496 93
rect 498 91 502 93
rect 493 83 502 91
rect 481 74 489 83
rect 481 72 484 74
rect 486 72 489 74
rect 481 70 489 72
rect 491 70 502 83
rect 504 83 509 95
rect 504 81 511 83
rect 504 79 507 81
rect 509 79 511 81
rect 530 80 535 95
rect 504 74 511 79
rect 504 72 507 74
rect 509 72 511 74
rect 504 70 511 72
rect 528 78 535 80
rect 528 76 530 78
rect 532 76 535 78
rect 528 71 535 76
rect 481 67 486 70
rect 528 69 530 71
rect 532 69 535 71
rect 528 67 535 69
rect 537 93 545 95
rect 537 91 540 93
rect 542 91 545 93
rect 537 86 545 91
rect 537 84 540 86
rect 542 84 545 86
rect 537 67 545 84
rect 547 85 555 95
rect 547 83 550 85
rect 552 83 555 85
rect 547 78 555 83
rect 547 76 550 78
rect 552 76 555 78
rect 547 67 555 76
rect 557 93 571 95
rect 557 91 562 93
rect 564 92 571 93
rect 594 93 603 95
rect 564 91 573 92
rect 557 86 573 91
rect 557 84 562 86
rect 564 84 573 86
rect 557 67 573 84
rect 575 67 580 92
rect 582 83 587 92
rect 594 91 597 93
rect 599 91 603 93
rect 594 83 603 91
rect 582 74 590 83
rect 582 72 585 74
rect 587 72 590 74
rect 582 70 590 72
rect 592 70 603 83
rect 605 83 610 95
rect 605 81 612 83
rect 605 79 608 81
rect 610 79 612 81
rect 629 80 634 95
rect 605 74 612 79
rect 605 72 608 74
rect 610 72 612 74
rect 605 70 612 72
rect 627 78 634 80
rect 627 76 629 78
rect 631 76 634 78
rect 627 71 634 76
rect 582 67 587 70
rect 627 69 629 71
rect 631 69 634 71
rect 627 67 634 69
rect 636 93 644 95
rect 636 91 639 93
rect 641 91 644 93
rect 636 86 644 91
rect 636 84 639 86
rect 641 84 644 86
rect 636 67 644 84
rect 646 85 654 95
rect 646 83 649 85
rect 651 83 654 85
rect 646 78 654 83
rect 646 76 649 78
rect 651 76 654 78
rect 646 67 654 76
rect 656 93 670 95
rect 656 91 661 93
rect 663 92 670 93
rect 693 93 702 95
rect 663 91 672 92
rect 656 86 672 91
rect 656 84 661 86
rect 663 84 672 86
rect 656 67 672 84
rect 674 67 679 92
rect 681 83 686 92
rect 693 91 696 93
rect 698 91 702 93
rect 693 83 702 91
rect 681 74 689 83
rect 681 72 684 74
rect 686 72 689 74
rect 681 70 689 72
rect 691 70 702 83
rect 704 83 709 95
rect 704 81 711 83
rect 704 79 707 81
rect 709 79 711 81
rect 704 74 711 79
rect 704 72 707 74
rect 709 72 711 74
rect 704 70 711 72
rect 681 67 686 70
<< alu1 >>
rect 362 390 366 391
rect 362 389 363 390
rect 27 388 363 389
rect 365 389 366 390
rect 408 390 412 391
rect 408 389 409 390
rect 365 388 409 389
rect 411 389 412 390
rect 453 390 457 391
rect 453 389 454 390
rect 411 388 454 389
rect 456 389 457 390
rect 526 390 530 391
rect 526 389 527 390
rect 456 388 527 389
rect 529 389 530 390
rect 529 388 716 389
rect 27 387 716 388
rect 27 386 68 387
rect 27 384 28 386
rect 30 385 68 386
rect 70 386 713 387
rect 70 385 106 386
rect 30 384 106 385
rect 108 384 177 386
rect 179 384 242 386
rect 244 384 295 386
rect 297 384 330 386
rect 332 384 592 386
rect 594 385 713 386
rect 715 385 716 387
rect 594 384 716 385
rect 27 381 716 384
rect 62 374 67 376
rect 62 372 63 374
rect 65 372 67 374
rect 31 359 35 368
rect 62 367 67 372
rect 102 374 107 376
rect 102 372 103 374
rect 105 372 107 374
rect 62 365 63 367
rect 65 365 67 367
rect 62 363 67 365
rect 31 358 44 359
rect 31 356 36 358
rect 38 356 41 358
rect 43 356 44 358
rect 31 355 44 356
rect 38 350 52 351
rect 38 348 46 350
rect 48 348 52 350
rect 38 347 52 348
rect 38 341 43 347
rect 38 339 39 341
rect 41 339 43 341
rect 38 338 43 339
rect 63 341 67 363
rect 71 359 75 368
rect 102 367 107 372
rect 183 371 196 375
rect 102 365 103 367
rect 105 365 107 367
rect 102 363 107 365
rect 71 358 84 359
rect 71 356 72 358
rect 74 356 76 358
rect 78 356 84 358
rect 71 355 84 356
rect 65 339 67 341
rect 63 336 67 339
rect 78 350 92 351
rect 78 348 86 350
rect 88 348 92 350
rect 78 347 92 348
rect 78 341 83 347
rect 78 339 79 341
rect 81 339 83 341
rect 78 338 83 339
rect 55 333 67 336
rect 103 341 107 363
rect 105 339 107 341
rect 103 336 107 339
rect 55 331 63 333
rect 65 331 67 333
rect 95 333 107 336
rect 95 331 103 333
rect 105 331 107 333
rect 111 366 117 368
rect 191 369 196 371
rect 191 367 192 369
rect 194 367 196 369
rect 111 364 114 366
rect 116 364 117 366
rect 111 359 117 364
rect 111 357 114 359
rect 116 357 117 359
rect 111 355 117 357
rect 111 335 115 355
rect 127 358 165 359
rect 127 356 128 358
rect 130 356 165 358
rect 127 355 165 356
rect 160 352 165 355
rect 135 350 150 351
rect 135 348 139 350
rect 141 348 146 350
rect 148 348 150 350
rect 135 347 150 348
rect 160 350 168 352
rect 160 348 165 350
rect 167 348 168 350
rect 144 341 148 347
rect 160 346 168 348
rect 191 362 196 367
rect 191 360 192 362
rect 194 360 196 362
rect 191 358 196 360
rect 144 339 145 341
rect 147 339 148 341
rect 144 338 148 339
rect 111 334 133 335
rect 111 332 114 334
rect 116 332 130 334
rect 132 332 133 334
rect 111 331 133 332
rect 192 336 196 358
rect 191 334 196 336
rect 191 332 192 334
rect 194 332 196 334
rect 55 330 67 331
rect 95 330 107 331
rect 191 330 196 332
rect 208 371 221 375
rect 297 374 302 376
rect 297 372 299 374
rect 301 372 302 374
rect 208 369 213 371
rect 208 367 210 369
rect 212 367 213 369
rect 208 362 213 367
rect 208 360 210 362
rect 212 360 213 362
rect 208 358 213 360
rect 208 336 212 358
rect 239 358 277 359
rect 239 356 274 358
rect 276 356 277 358
rect 239 355 277 356
rect 239 352 244 355
rect 236 350 244 352
rect 236 348 237 350
rect 239 348 244 350
rect 236 346 244 348
rect 254 350 269 351
rect 254 348 256 350
rect 258 348 263 350
rect 265 348 269 350
rect 254 347 269 348
rect 208 334 213 336
rect 256 341 260 347
rect 287 366 293 368
rect 287 364 288 366
rect 290 364 293 366
rect 287 359 293 364
rect 287 357 288 359
rect 290 357 293 359
rect 287 355 293 357
rect 256 339 257 341
rect 259 339 260 341
rect 256 338 260 339
rect 289 335 293 355
rect 208 332 210 334
rect 212 332 213 334
rect 208 330 213 332
rect 271 334 293 335
rect 271 332 272 334
rect 274 332 288 334
rect 290 332 293 334
rect 271 331 293 332
rect 297 367 302 372
rect 337 374 342 376
rect 337 372 339 374
rect 341 372 342 374
rect 297 365 299 367
rect 301 365 302 367
rect 297 363 302 365
rect 297 341 301 363
rect 329 359 333 368
rect 320 358 333 359
rect 320 356 326 358
rect 328 356 330 358
rect 332 356 333 358
rect 320 355 333 356
rect 337 367 342 372
rect 378 371 391 375
rect 467 374 472 376
rect 467 372 469 374
rect 471 372 472 374
rect 378 369 383 371
rect 337 365 339 367
rect 341 365 342 367
rect 337 363 342 365
rect 312 350 326 351
rect 312 348 316 350
rect 318 348 326 350
rect 312 347 326 348
rect 297 339 299 341
rect 297 336 301 339
rect 297 333 309 336
rect 297 331 299 333
rect 301 331 309 333
rect 321 341 326 347
rect 321 339 323 341
rect 325 339 326 341
rect 321 338 326 339
rect 337 341 341 363
rect 369 359 373 368
rect 360 358 373 359
rect 360 356 361 358
rect 363 356 366 358
rect 368 356 373 358
rect 360 355 373 356
rect 378 367 380 369
rect 382 367 383 369
rect 378 362 383 367
rect 378 360 380 362
rect 382 360 383 362
rect 378 358 383 360
rect 352 350 366 351
rect 352 348 356 350
rect 358 348 366 350
rect 352 347 366 348
rect 337 339 339 341
rect 337 336 341 339
rect 337 333 349 336
rect 337 331 339 333
rect 341 331 349 333
rect 361 341 366 347
rect 361 339 363 341
rect 365 339 366 341
rect 361 338 366 339
rect 378 336 382 358
rect 409 358 447 359
rect 409 356 444 358
rect 446 356 447 358
rect 409 355 447 356
rect 409 352 414 355
rect 406 350 414 352
rect 406 348 407 350
rect 409 348 414 350
rect 406 346 414 348
rect 424 350 439 351
rect 424 348 426 350
rect 428 348 433 350
rect 435 348 439 350
rect 424 347 439 348
rect 378 334 383 336
rect 426 341 430 347
rect 457 366 463 368
rect 457 364 458 366
rect 460 364 463 366
rect 457 359 463 364
rect 457 357 458 359
rect 460 357 463 359
rect 457 355 463 357
rect 426 339 427 341
rect 429 339 430 341
rect 426 338 430 339
rect 459 335 463 355
rect 378 332 380 334
rect 382 332 383 334
rect 297 330 309 331
rect 337 330 349 331
rect 378 330 383 332
rect 441 334 463 335
rect 441 332 442 334
rect 444 332 458 334
rect 460 332 463 334
rect 441 331 463 332
rect 467 367 472 372
rect 507 374 512 376
rect 507 372 509 374
rect 511 372 512 374
rect 467 365 469 367
rect 471 365 472 367
rect 467 363 472 365
rect 467 341 471 363
rect 499 359 503 368
rect 490 358 503 359
rect 490 356 496 358
rect 498 356 500 358
rect 502 356 503 358
rect 490 355 503 356
rect 507 367 512 372
rect 578 374 583 376
rect 578 372 579 374
rect 581 372 583 374
rect 507 365 509 367
rect 511 365 512 367
rect 507 363 512 365
rect 482 350 496 351
rect 482 348 486 350
rect 488 348 496 350
rect 482 347 496 348
rect 467 339 469 341
rect 467 336 471 339
rect 467 333 479 336
rect 467 331 469 333
rect 471 331 479 333
rect 491 341 496 347
rect 491 339 493 341
rect 495 339 496 341
rect 491 338 496 339
rect 507 341 511 363
rect 539 359 543 368
rect 530 358 543 359
rect 530 356 531 358
rect 533 356 536 358
rect 538 356 543 358
rect 530 355 543 356
rect 547 359 551 368
rect 578 367 583 372
rect 618 374 623 376
rect 618 372 619 374
rect 621 372 623 374
rect 578 365 579 367
rect 581 365 583 367
rect 578 363 583 365
rect 547 358 560 359
rect 547 356 552 358
rect 554 356 557 358
rect 559 356 560 358
rect 547 355 560 356
rect 522 350 536 351
rect 522 348 526 350
rect 528 348 536 350
rect 522 347 536 348
rect 507 339 509 341
rect 507 336 511 339
rect 507 333 519 336
rect 507 331 509 333
rect 511 331 519 333
rect 531 341 536 347
rect 531 339 533 341
rect 535 339 536 341
rect 531 338 536 339
rect 554 350 568 351
rect 554 348 562 350
rect 564 348 568 350
rect 554 347 568 348
rect 554 341 559 347
rect 554 339 555 341
rect 557 339 559 341
rect 554 338 559 339
rect 579 341 583 363
rect 587 359 591 368
rect 618 367 623 372
rect 699 371 712 375
rect 618 365 619 367
rect 621 365 623 367
rect 618 363 623 365
rect 587 358 600 359
rect 587 356 588 358
rect 590 356 592 358
rect 594 356 600 358
rect 587 355 600 356
rect 581 339 583 341
rect 579 336 583 339
rect 594 350 608 351
rect 594 348 602 350
rect 604 348 608 350
rect 594 347 608 348
rect 594 341 599 347
rect 594 339 595 341
rect 597 339 599 341
rect 594 338 599 339
rect 571 333 583 336
rect 619 341 623 363
rect 621 339 623 341
rect 619 336 623 339
rect 571 331 579 333
rect 581 331 583 333
rect 611 333 623 336
rect 611 331 619 333
rect 621 331 623 333
rect 627 366 633 368
rect 707 369 712 371
rect 707 367 708 369
rect 710 367 712 369
rect 627 364 630 366
rect 632 364 633 366
rect 627 359 633 364
rect 627 357 630 359
rect 632 357 633 359
rect 627 355 633 357
rect 627 335 631 355
rect 643 358 681 359
rect 643 356 644 358
rect 646 356 681 358
rect 643 355 681 356
rect 676 352 681 355
rect 651 350 666 351
rect 651 348 655 350
rect 657 348 662 350
rect 664 348 666 350
rect 651 347 666 348
rect 676 350 684 352
rect 676 348 681 350
rect 683 348 684 350
rect 660 341 664 347
rect 676 346 684 348
rect 707 362 712 367
rect 707 360 708 362
rect 710 360 712 362
rect 707 358 712 360
rect 660 339 661 341
rect 663 339 664 341
rect 660 338 664 339
rect 627 334 649 335
rect 627 332 630 334
rect 632 332 646 334
rect 648 332 649 334
rect 627 331 649 332
rect 708 336 712 358
rect 707 334 712 336
rect 707 332 708 334
rect 710 332 712 334
rect 467 330 479 331
rect 507 330 519 331
rect 571 330 583 331
rect 611 330 623 331
rect 707 330 712 332
rect 27 324 716 325
rect 27 322 52 324
rect 54 322 92 324
rect 94 322 310 324
rect 312 322 350 324
rect 352 322 480 324
rect 482 322 520 324
rect 522 322 568 324
rect 570 322 608 324
rect 610 322 716 324
rect 27 318 716 322
rect 27 316 28 318
rect 30 316 89 318
rect 91 316 153 318
rect 155 316 217 318
rect 219 316 280 318
rect 282 316 315 318
rect 317 316 347 318
rect 349 316 388 318
rect 390 316 419 318
rect 421 316 476 318
rect 478 316 566 318
rect 568 316 669 318
rect 671 316 713 318
rect 715 316 716 318
rect 27 312 716 316
rect 27 310 52 312
rect 54 310 92 312
rect 94 310 310 312
rect 312 310 350 312
rect 352 310 480 312
rect 482 310 520 312
rect 522 310 568 312
rect 570 310 608 312
rect 610 310 716 312
rect 27 309 716 310
rect 55 303 67 304
rect 95 303 107 304
rect 38 295 43 296
rect 38 293 39 295
rect 41 293 43 295
rect 38 287 43 293
rect 55 301 63 303
rect 65 301 67 303
rect 55 298 67 301
rect 63 295 67 298
rect 65 293 67 295
rect 38 286 52 287
rect 38 284 46 286
rect 48 284 52 286
rect 38 283 52 284
rect 31 278 44 279
rect 31 276 36 278
rect 38 276 41 278
rect 43 276 44 278
rect 31 275 44 276
rect 63 286 67 293
rect 63 284 64 286
rect 66 284 67 286
rect 31 266 35 275
rect 63 271 67 284
rect 78 295 83 296
rect 78 293 79 295
rect 81 293 83 295
rect 78 287 83 293
rect 95 301 103 303
rect 105 301 107 303
rect 95 298 107 301
rect 103 295 107 298
rect 105 293 107 295
rect 78 286 92 287
rect 78 284 86 286
rect 88 284 92 286
rect 78 283 92 284
rect 62 269 67 271
rect 62 267 63 269
rect 65 267 67 269
rect 62 262 67 267
rect 71 278 84 279
rect 71 276 72 278
rect 74 276 76 278
rect 78 276 84 278
rect 71 275 84 276
rect 71 266 75 275
rect 103 271 107 293
rect 102 269 107 271
rect 102 267 103 269
rect 105 267 107 269
rect 62 260 63 262
rect 65 260 67 262
rect 62 258 67 260
rect 102 262 107 267
rect 111 302 133 303
rect 111 300 114 302
rect 116 300 133 302
rect 111 299 133 300
rect 191 302 196 304
rect 191 300 192 302
rect 194 300 196 302
rect 111 279 115 299
rect 111 277 117 279
rect 111 275 114 277
rect 116 275 117 277
rect 111 270 117 275
rect 111 268 114 270
rect 116 268 117 270
rect 111 266 117 268
rect 144 287 148 296
rect 191 298 196 300
rect 135 286 150 287
rect 135 284 136 286
rect 138 284 139 286
rect 141 284 146 286
rect 148 284 150 286
rect 135 283 150 284
rect 160 286 168 288
rect 160 284 165 286
rect 167 284 168 286
rect 160 282 168 284
rect 160 279 165 282
rect 127 278 165 279
rect 127 276 128 278
rect 130 276 165 278
rect 127 275 165 276
rect 192 276 196 298
rect 191 274 196 276
rect 191 272 192 274
rect 194 272 196 274
rect 191 267 196 272
rect 191 265 192 267
rect 194 265 196 267
rect 191 263 196 265
rect 102 260 103 262
rect 105 260 107 262
rect 102 258 107 260
rect 183 259 196 263
rect 208 302 213 304
rect 297 303 309 304
rect 337 303 349 304
rect 208 300 210 302
rect 212 300 213 302
rect 208 298 213 300
rect 208 276 212 298
rect 271 302 293 303
rect 271 300 288 302
rect 290 300 293 302
rect 271 299 293 300
rect 208 274 213 276
rect 208 272 210 274
rect 212 272 213 274
rect 208 267 213 272
rect 236 286 244 288
rect 256 287 260 296
rect 236 284 237 286
rect 239 284 244 286
rect 236 282 244 284
rect 254 286 269 287
rect 254 284 256 286
rect 258 284 263 286
rect 265 284 266 286
rect 268 284 269 286
rect 254 283 269 284
rect 239 279 244 282
rect 239 278 277 279
rect 239 276 274 278
rect 276 276 277 278
rect 239 275 277 276
rect 289 279 293 299
rect 287 277 293 279
rect 287 275 288 277
rect 290 275 293 277
rect 287 270 293 275
rect 287 268 288 270
rect 290 268 293 270
rect 208 265 210 267
rect 212 265 213 267
rect 208 263 213 265
rect 287 266 293 268
rect 297 301 299 303
rect 301 301 309 303
rect 297 298 309 301
rect 337 301 339 303
rect 341 301 349 303
rect 297 295 301 298
rect 297 293 299 295
rect 297 271 301 293
rect 337 298 349 301
rect 378 302 383 304
rect 467 303 479 304
rect 507 303 519 304
rect 571 303 583 304
rect 611 303 623 304
rect 378 300 380 302
rect 382 300 383 302
rect 321 295 326 296
rect 321 293 323 295
rect 325 293 326 295
rect 321 287 326 293
rect 312 286 326 287
rect 312 284 316 286
rect 318 284 326 286
rect 312 283 326 284
rect 337 295 341 298
rect 337 293 339 295
rect 320 278 333 279
rect 320 276 326 278
rect 328 276 330 278
rect 332 276 333 278
rect 320 275 333 276
rect 297 269 302 271
rect 297 267 299 269
rect 301 267 302 269
rect 208 259 221 263
rect 297 262 302 267
rect 329 266 333 275
rect 337 271 341 293
rect 378 298 383 300
rect 361 295 366 296
rect 361 293 363 295
rect 365 293 366 295
rect 361 287 366 293
rect 352 286 366 287
rect 352 284 356 286
rect 358 284 366 286
rect 352 283 366 284
rect 360 278 373 279
rect 360 276 361 278
rect 363 276 366 278
rect 368 276 373 278
rect 360 275 373 276
rect 337 269 342 271
rect 337 267 339 269
rect 341 267 342 269
rect 297 260 299 262
rect 301 260 302 262
rect 297 258 302 260
rect 337 265 342 267
rect 337 263 339 265
rect 341 263 342 265
rect 369 266 373 275
rect 378 276 382 298
rect 441 302 463 303
rect 441 300 458 302
rect 460 300 463 302
rect 441 299 463 300
rect 378 274 383 276
rect 378 272 380 274
rect 382 272 383 274
rect 378 267 383 272
rect 406 286 414 288
rect 426 287 430 296
rect 459 294 463 299
rect 459 292 460 294
rect 462 292 463 294
rect 406 284 407 286
rect 409 284 414 286
rect 406 282 414 284
rect 424 286 439 287
rect 424 284 426 286
rect 428 284 433 286
rect 435 284 436 286
rect 438 284 439 286
rect 424 283 439 284
rect 409 279 414 282
rect 409 278 447 279
rect 409 276 444 278
rect 446 276 447 278
rect 409 275 447 276
rect 459 279 463 292
rect 457 277 463 279
rect 457 275 458 277
rect 460 275 463 277
rect 457 270 463 275
rect 457 268 458 270
rect 460 268 463 270
rect 337 262 342 263
rect 337 260 339 262
rect 341 260 342 262
rect 337 258 342 260
rect 378 265 380 267
rect 382 265 383 267
rect 378 263 383 265
rect 457 266 463 268
rect 467 301 469 303
rect 471 301 479 303
rect 467 298 479 301
rect 507 301 509 303
rect 511 301 519 303
rect 467 295 471 298
rect 467 293 469 295
rect 467 271 471 293
rect 507 298 519 301
rect 491 295 496 296
rect 491 293 493 295
rect 495 293 496 295
rect 491 287 496 293
rect 482 286 496 287
rect 482 284 486 286
rect 488 284 496 286
rect 482 283 496 284
rect 507 295 511 298
rect 507 293 509 295
rect 507 286 511 293
rect 531 295 536 296
rect 531 293 533 295
rect 535 293 536 295
rect 507 284 508 286
rect 510 284 511 286
rect 490 278 503 279
rect 490 276 496 278
rect 498 276 500 278
rect 502 276 503 278
rect 490 275 503 276
rect 467 269 472 271
rect 467 267 469 269
rect 471 267 472 269
rect 378 259 391 263
rect 467 262 472 267
rect 499 266 503 275
rect 507 271 511 284
rect 531 287 536 293
rect 522 286 536 287
rect 522 284 526 286
rect 528 284 536 286
rect 522 283 536 284
rect 554 295 559 296
rect 554 293 555 295
rect 557 293 559 295
rect 554 287 559 293
rect 571 301 579 303
rect 581 301 583 303
rect 571 298 583 301
rect 579 295 583 298
rect 581 293 583 295
rect 554 286 568 287
rect 554 284 562 286
rect 564 284 568 286
rect 554 283 568 284
rect 530 278 543 279
rect 530 276 531 278
rect 533 276 536 278
rect 538 276 543 278
rect 530 275 543 276
rect 507 269 512 271
rect 507 267 509 269
rect 511 267 512 269
rect 467 260 469 262
rect 471 260 472 262
rect 467 258 472 260
rect 507 262 512 267
rect 539 266 543 275
rect 547 278 560 279
rect 547 276 552 278
rect 554 276 557 278
rect 559 276 560 278
rect 547 275 560 276
rect 547 266 551 275
rect 579 271 583 293
rect 594 295 599 296
rect 594 293 595 295
rect 597 293 599 295
rect 594 287 599 293
rect 611 301 619 303
rect 621 301 623 303
rect 611 298 623 301
rect 619 295 623 298
rect 621 293 623 295
rect 594 286 608 287
rect 594 284 602 286
rect 604 284 608 286
rect 594 283 608 284
rect 578 269 583 271
rect 578 267 579 269
rect 581 267 583 269
rect 507 260 509 262
rect 511 260 512 262
rect 507 258 512 260
rect 578 262 583 267
rect 587 278 600 279
rect 587 276 588 278
rect 590 276 592 278
rect 594 276 600 278
rect 587 275 600 276
rect 587 266 591 275
rect 619 271 623 293
rect 618 269 623 271
rect 618 267 619 269
rect 621 267 623 269
rect 578 260 579 262
rect 581 260 583 262
rect 578 258 583 260
rect 618 262 623 267
rect 627 302 649 303
rect 627 300 630 302
rect 632 300 649 302
rect 627 299 649 300
rect 707 302 712 304
rect 707 300 708 302
rect 710 300 712 302
rect 627 279 631 299
rect 627 277 633 279
rect 627 275 630 277
rect 632 275 633 277
rect 627 270 633 275
rect 627 268 630 270
rect 632 268 633 270
rect 627 266 633 268
rect 660 287 664 296
rect 707 298 712 300
rect 651 286 666 287
rect 651 284 652 286
rect 654 284 655 286
rect 657 284 662 286
rect 664 284 666 286
rect 651 283 666 284
rect 676 286 684 288
rect 676 284 681 286
rect 683 284 684 286
rect 676 282 684 284
rect 676 279 681 282
rect 643 278 681 279
rect 643 276 644 278
rect 646 276 681 278
rect 643 275 681 276
rect 708 276 712 298
rect 707 274 712 276
rect 707 272 708 274
rect 710 272 712 274
rect 707 267 712 272
rect 707 265 708 267
rect 710 265 712 267
rect 707 263 712 265
rect 618 260 619 262
rect 621 260 623 262
rect 618 258 623 260
rect 699 262 712 263
rect 699 260 700 262
rect 702 260 712 262
rect 699 259 712 260
rect 27 247 716 253
rect 27 246 713 247
rect 27 245 68 246
rect 27 243 28 245
rect 30 244 68 245
rect 70 244 106 246
rect 108 244 177 246
rect 179 244 242 246
rect 244 244 295 246
rect 297 245 409 246
rect 297 244 330 245
rect 30 243 330 244
rect 332 243 362 245
rect 364 244 409 245
rect 411 244 454 246
rect 456 245 713 246
rect 715 245 716 247
rect 456 244 527 245
rect 364 243 527 244
rect 529 243 592 245
rect 594 243 716 245
rect 27 240 716 243
rect 27 238 44 240
rect 46 238 388 240
rect 390 238 716 240
rect 27 237 716 238
rect 31 231 43 232
rect 31 229 33 231
rect 35 229 43 231
rect 31 226 43 229
rect 31 224 35 226
rect 31 222 33 224
rect 31 199 35 222
rect 143 230 156 231
rect 143 228 153 230
rect 155 228 156 230
rect 143 227 156 228
rect 244 227 257 231
rect 375 231 387 232
rect 346 227 359 231
rect 55 222 77 224
rect 151 225 156 227
rect 151 223 152 225
rect 154 223 156 225
rect 55 220 74 222
rect 76 220 77 222
rect 55 218 67 220
rect 31 197 36 199
rect 31 195 33 197
rect 35 195 36 197
rect 31 190 36 195
rect 47 208 51 216
rect 47 206 59 208
rect 47 204 50 206
rect 52 205 59 206
rect 52 204 53 205
rect 47 203 53 204
rect 55 203 59 205
rect 47 202 59 203
rect 63 206 67 218
rect 65 204 67 206
rect 63 202 67 204
rect 71 215 77 220
rect 71 213 74 215
rect 76 213 77 215
rect 71 211 77 213
rect 31 188 33 190
rect 35 188 36 190
rect 31 186 36 188
rect 71 191 75 211
rect 87 214 125 215
rect 87 212 122 214
rect 124 212 125 214
rect 87 211 125 212
rect 120 208 125 211
rect 95 206 110 207
rect 95 204 99 206
rect 101 204 106 206
rect 108 204 110 206
rect 95 203 110 204
rect 120 206 128 208
rect 120 204 125 206
rect 127 204 128 206
rect 104 197 108 203
rect 120 202 128 204
rect 151 218 156 223
rect 151 216 152 218
rect 154 216 156 218
rect 151 214 156 216
rect 104 195 105 197
rect 107 195 108 197
rect 104 194 108 195
rect 71 190 93 191
rect 71 188 74 190
rect 76 188 93 190
rect 71 187 93 188
rect 152 192 156 214
rect 151 190 156 192
rect 151 188 152 190
rect 154 188 156 190
rect 151 186 156 188
rect 172 222 178 224
rect 252 225 257 227
rect 252 223 253 225
rect 255 223 257 225
rect 172 220 175 222
rect 177 220 178 222
rect 172 215 178 220
rect 172 213 175 215
rect 177 213 178 215
rect 172 211 178 213
rect 172 191 176 211
rect 188 214 226 215
rect 188 212 210 214
rect 212 212 226 214
rect 188 211 226 212
rect 221 208 226 211
rect 196 206 211 207
rect 196 204 200 206
rect 202 204 207 206
rect 209 204 211 206
rect 196 203 211 204
rect 221 206 229 208
rect 221 204 226 206
rect 228 204 229 206
rect 205 194 209 203
rect 221 202 229 204
rect 252 218 257 223
rect 252 216 253 218
rect 255 216 257 218
rect 252 214 257 216
rect 172 190 194 191
rect 172 188 175 190
rect 177 188 194 190
rect 172 187 194 188
rect 253 192 257 214
rect 252 190 257 192
rect 252 188 253 190
rect 255 188 257 190
rect 252 186 257 188
rect 274 222 280 224
rect 354 225 359 227
rect 354 223 355 225
rect 357 223 359 225
rect 274 220 277 222
rect 279 220 280 222
rect 274 215 280 220
rect 274 213 277 215
rect 279 213 280 215
rect 274 211 280 213
rect 274 191 278 211
rect 290 214 328 215
rect 290 212 291 214
rect 293 212 328 214
rect 290 211 328 212
rect 323 208 328 211
rect 298 206 313 207
rect 298 204 302 206
rect 304 204 309 206
rect 311 204 313 206
rect 298 203 313 204
rect 323 206 331 208
rect 323 204 328 206
rect 330 204 331 206
rect 307 197 311 203
rect 323 202 331 204
rect 354 218 359 223
rect 354 216 355 218
rect 357 216 359 218
rect 354 214 359 216
rect 307 195 308 197
rect 310 195 311 197
rect 307 194 311 195
rect 274 190 296 191
rect 274 188 277 190
rect 279 188 296 190
rect 274 187 296 188
rect 355 192 359 214
rect 354 190 359 192
rect 354 188 355 190
rect 357 188 359 190
rect 354 186 359 188
rect 375 229 377 231
rect 379 229 387 231
rect 375 226 387 229
rect 375 224 379 226
rect 375 222 377 224
rect 375 206 379 222
rect 499 227 512 231
rect 600 227 613 231
rect 699 227 712 231
rect 375 204 376 206
rect 378 204 379 206
rect 375 199 379 204
rect 399 222 433 224
rect 507 225 512 227
rect 507 223 508 225
rect 510 223 512 225
rect 399 220 430 222
rect 432 220 433 222
rect 399 218 411 220
rect 375 197 380 199
rect 375 195 377 197
rect 379 195 380 197
rect 375 190 380 195
rect 391 208 395 216
rect 391 206 403 208
rect 391 204 394 206
rect 396 205 403 206
rect 396 204 399 205
rect 391 203 399 204
rect 401 203 403 205
rect 391 202 403 203
rect 407 206 411 218
rect 409 204 411 206
rect 407 202 411 204
rect 427 215 433 220
rect 427 213 430 215
rect 432 213 433 215
rect 427 211 433 213
rect 375 188 377 190
rect 379 188 380 190
rect 375 186 380 188
rect 427 191 431 211
rect 443 214 481 215
rect 443 212 444 214
rect 446 212 481 214
rect 443 211 481 212
rect 476 208 481 211
rect 451 206 466 207
rect 451 204 455 206
rect 457 204 462 206
rect 464 204 466 206
rect 451 203 466 204
rect 476 206 484 208
rect 476 204 481 206
rect 483 204 484 206
rect 460 194 464 203
rect 476 202 484 204
rect 507 218 512 223
rect 507 216 508 218
rect 510 216 512 218
rect 507 214 512 216
rect 427 190 449 191
rect 427 188 430 190
rect 432 188 449 190
rect 427 187 449 188
rect 508 192 512 214
rect 507 190 512 192
rect 504 189 508 190
rect 504 187 505 189
rect 507 188 508 189
rect 510 188 512 190
rect 507 187 512 188
rect 528 222 534 224
rect 608 225 613 227
rect 608 223 609 225
rect 611 223 613 225
rect 528 220 531 222
rect 533 220 534 222
rect 528 215 534 220
rect 528 213 531 215
rect 533 213 534 215
rect 528 211 534 213
rect 528 197 532 211
rect 544 214 582 215
rect 544 212 545 214
rect 547 212 582 214
rect 544 211 582 212
rect 577 208 582 211
rect 552 206 567 207
rect 552 204 556 206
rect 558 204 563 206
rect 565 204 567 206
rect 552 203 567 204
rect 577 206 585 208
rect 577 204 582 206
rect 584 204 585 206
rect 528 195 529 197
rect 531 195 532 197
rect 528 191 532 195
rect 561 197 565 203
rect 577 202 585 204
rect 608 218 613 223
rect 608 216 609 218
rect 611 216 613 218
rect 608 214 613 216
rect 609 205 613 214
rect 609 203 610 205
rect 612 203 613 205
rect 561 195 562 197
rect 564 195 565 197
rect 561 194 565 195
rect 528 190 550 191
rect 528 188 531 190
rect 533 188 550 190
rect 528 187 550 188
rect 609 192 613 203
rect 608 190 613 192
rect 608 188 609 190
rect 611 188 613 190
rect 504 186 512 187
rect 608 186 613 188
rect 627 222 633 224
rect 707 225 712 227
rect 707 223 708 225
rect 710 223 712 225
rect 627 220 630 222
rect 632 220 633 222
rect 627 215 633 220
rect 627 213 630 215
rect 632 213 633 215
rect 627 211 633 213
rect 627 197 631 211
rect 643 214 681 215
rect 643 212 644 214
rect 646 212 681 214
rect 643 211 681 212
rect 676 208 681 211
rect 651 206 666 207
rect 651 204 652 206
rect 654 204 655 206
rect 657 204 662 206
rect 664 204 666 206
rect 651 203 666 204
rect 676 206 684 208
rect 676 204 681 206
rect 683 204 684 206
rect 627 195 628 197
rect 630 195 631 197
rect 627 191 631 195
rect 660 194 664 203
rect 676 202 684 204
rect 707 218 712 223
rect 707 216 708 218
rect 710 216 712 218
rect 707 214 712 216
rect 627 190 649 191
rect 627 188 630 190
rect 632 188 649 190
rect 627 187 649 188
rect 708 192 712 214
rect 707 190 712 192
rect 707 188 708 190
rect 710 188 712 190
rect 707 186 712 188
rect 27 180 716 181
rect 27 178 404 180
rect 406 178 716 180
rect 27 175 716 178
rect 24 174 716 175
rect 24 172 25 174
rect 27 173 153 174
rect 27 172 89 173
rect 24 171 89 172
rect 91 172 153 173
rect 155 172 217 174
rect 219 172 280 174
rect 282 172 316 174
rect 318 172 347 174
rect 349 173 566 174
rect 349 172 388 173
rect 91 171 388 172
rect 390 171 419 173
rect 421 171 476 173
rect 478 172 566 173
rect 568 172 669 174
rect 671 172 713 174
rect 715 172 716 174
rect 478 171 716 172
rect 27 168 716 171
rect 27 166 150 168
rect 152 166 404 168
rect 406 166 716 168
rect 27 165 716 166
rect 32 158 54 159
rect 32 156 35 158
rect 37 156 51 158
rect 53 156 54 158
rect 32 155 54 156
rect 112 158 117 160
rect 112 156 113 158
rect 115 156 117 158
rect 32 135 36 155
rect 65 150 69 152
rect 65 148 66 150
rect 68 148 69 150
rect 32 133 38 135
rect 32 131 35 133
rect 37 131 38 133
rect 32 126 38 131
rect 32 124 35 126
rect 37 124 38 126
rect 32 122 38 124
rect 65 143 69 148
rect 112 154 117 156
rect 56 142 71 143
rect 56 140 60 142
rect 62 140 67 142
rect 69 140 71 142
rect 56 139 71 140
rect 81 142 89 144
rect 81 140 86 142
rect 88 140 89 142
rect 81 138 89 140
rect 81 135 86 138
rect 48 134 86 135
rect 48 132 83 134
rect 85 132 86 134
rect 48 131 86 132
rect 113 132 117 154
rect 112 130 117 132
rect 112 128 113 130
rect 115 128 117 130
rect 112 123 117 128
rect 112 121 113 123
rect 115 121 117 123
rect 112 119 117 121
rect 104 115 117 119
rect 121 158 126 160
rect 121 156 123 158
rect 125 156 126 158
rect 121 151 126 156
rect 173 158 195 159
rect 173 156 176 158
rect 178 156 195 158
rect 173 155 195 156
rect 253 158 258 160
rect 253 156 254 158
rect 256 156 258 158
rect 121 149 123 151
rect 125 149 126 151
rect 121 147 126 149
rect 121 124 125 147
rect 173 144 177 155
rect 206 151 210 152
rect 206 149 207 151
rect 209 149 210 151
rect 137 143 149 144
rect 137 142 145 143
rect 137 140 140 142
rect 142 141 145 142
rect 147 141 149 143
rect 142 140 149 141
rect 137 138 149 140
rect 137 130 141 138
rect 153 142 177 144
rect 155 140 177 142
rect 153 128 157 140
rect 121 122 123 124
rect 121 120 125 122
rect 121 117 133 120
rect 121 115 123 117
rect 125 115 133 117
rect 121 114 133 115
rect 145 122 157 128
rect 173 135 177 140
rect 173 133 179 135
rect 173 131 176 133
rect 178 131 179 133
rect 173 126 179 131
rect 173 124 176 126
rect 178 124 179 126
rect 173 122 179 124
rect 206 143 210 149
rect 253 154 258 156
rect 254 150 258 154
rect 254 148 255 150
rect 257 148 258 150
rect 197 142 212 143
rect 197 140 201 142
rect 203 140 208 142
rect 210 140 212 142
rect 197 139 212 140
rect 222 142 230 144
rect 222 140 227 142
rect 229 140 230 142
rect 222 138 230 140
rect 222 135 227 138
rect 189 131 227 135
rect 254 132 258 148
rect 253 130 258 132
rect 253 128 254 130
rect 256 128 258 130
rect 253 123 258 128
rect 253 121 254 123
rect 256 121 258 123
rect 253 119 258 121
rect 245 115 258 119
rect 274 158 279 160
rect 274 156 276 158
rect 278 156 279 158
rect 274 154 279 156
rect 274 132 278 154
rect 337 158 359 159
rect 337 156 338 158
rect 340 156 354 158
rect 356 156 359 158
rect 337 155 359 156
rect 322 150 326 152
rect 322 148 323 150
rect 325 148 326 150
rect 274 130 279 132
rect 274 128 276 130
rect 278 128 279 130
rect 274 123 279 128
rect 302 142 310 144
rect 322 143 326 148
rect 302 140 303 142
rect 305 140 310 142
rect 302 138 310 140
rect 320 142 335 143
rect 320 140 322 142
rect 324 140 329 142
rect 331 140 335 142
rect 320 139 335 140
rect 305 135 310 138
rect 305 134 343 135
rect 305 132 340 134
rect 342 132 343 134
rect 305 131 343 132
rect 355 135 359 155
rect 353 133 359 135
rect 353 131 354 133
rect 356 131 359 133
rect 353 126 359 131
rect 353 124 354 126
rect 356 124 359 126
rect 274 121 276 123
rect 278 121 279 123
rect 274 119 279 121
rect 353 122 359 124
rect 375 158 380 160
rect 375 156 377 158
rect 379 156 380 158
rect 375 151 380 156
rect 427 158 449 159
rect 427 156 430 158
rect 432 156 449 158
rect 427 155 449 156
rect 507 158 512 160
rect 507 156 508 158
rect 510 156 512 158
rect 375 149 377 151
rect 379 149 380 151
rect 375 147 380 149
rect 375 134 379 147
rect 375 132 376 134
rect 378 132 379 134
rect 375 124 379 132
rect 391 143 403 144
rect 391 142 399 143
rect 391 140 394 142
rect 396 141 399 142
rect 401 141 403 143
rect 396 140 403 141
rect 391 138 403 140
rect 391 130 395 138
rect 407 142 411 144
rect 409 140 411 142
rect 407 128 411 140
rect 375 122 377 124
rect 375 120 379 122
rect 274 118 287 119
rect 274 116 284 118
rect 286 116 287 118
rect 274 115 287 116
rect 375 117 387 120
rect 375 115 377 117
rect 379 115 387 117
rect 375 114 387 115
rect 399 126 411 128
rect 427 135 431 155
rect 427 133 433 135
rect 427 131 430 133
rect 432 131 433 133
rect 427 126 433 131
rect 399 124 430 126
rect 432 124 433 126
rect 399 122 433 124
rect 460 143 464 152
rect 507 154 512 156
rect 451 142 466 143
rect 451 140 455 142
rect 457 140 462 142
rect 464 140 466 142
rect 451 139 466 140
rect 476 142 484 144
rect 476 140 481 142
rect 483 140 484 142
rect 476 138 484 140
rect 476 135 481 138
rect 443 134 481 135
rect 443 132 478 134
rect 480 132 481 134
rect 443 131 481 132
rect 508 132 512 154
rect 507 130 512 132
rect 507 128 508 130
rect 510 128 512 130
rect 507 123 512 128
rect 507 121 508 123
rect 510 121 512 123
rect 528 158 550 159
rect 528 156 531 158
rect 533 156 550 158
rect 528 155 550 156
rect 608 158 613 160
rect 608 156 609 158
rect 611 156 613 158
rect 528 151 532 155
rect 528 149 529 151
rect 531 149 532 151
rect 528 135 532 149
rect 561 151 565 152
rect 561 149 562 151
rect 564 149 565 151
rect 528 133 534 135
rect 528 131 531 133
rect 533 131 534 133
rect 528 126 534 131
rect 528 124 531 126
rect 533 124 534 126
rect 528 122 534 124
rect 561 143 565 149
rect 608 154 613 156
rect 552 142 567 143
rect 552 140 556 142
rect 558 140 563 142
rect 565 140 567 142
rect 552 139 567 140
rect 577 142 585 144
rect 577 140 582 142
rect 584 140 585 142
rect 577 138 585 140
rect 577 135 582 138
rect 609 143 613 154
rect 609 141 610 143
rect 612 141 613 143
rect 544 133 579 135
rect 581 133 582 135
rect 544 131 582 133
rect 609 132 613 141
rect 608 130 613 132
rect 608 128 609 130
rect 611 128 613 130
rect 608 123 613 128
rect 507 119 512 121
rect 608 121 609 123
rect 611 121 613 123
rect 627 158 649 159
rect 627 156 630 158
rect 632 156 649 158
rect 627 155 649 156
rect 707 158 712 160
rect 707 156 708 158
rect 710 156 712 158
rect 627 151 631 155
rect 627 149 628 151
rect 630 149 631 151
rect 627 135 631 149
rect 660 151 664 152
rect 660 149 661 151
rect 663 149 664 151
rect 627 133 633 135
rect 627 131 630 133
rect 632 131 633 133
rect 627 126 633 131
rect 627 124 630 126
rect 632 124 633 126
rect 627 122 633 124
rect 660 143 664 149
rect 707 154 712 156
rect 651 142 666 143
rect 651 140 655 142
rect 657 140 662 142
rect 664 140 666 142
rect 651 139 666 140
rect 676 142 684 144
rect 676 140 681 142
rect 683 140 684 142
rect 676 138 684 140
rect 676 135 681 138
rect 643 134 681 135
rect 643 132 678 134
rect 680 132 681 134
rect 643 131 681 132
rect 708 132 712 154
rect 707 130 712 132
rect 707 128 708 130
rect 710 128 712 130
rect 707 123 712 128
rect 608 119 613 121
rect 707 121 708 123
rect 710 121 712 123
rect 707 119 712 121
rect 499 115 512 119
rect 600 115 613 119
rect 699 115 712 119
rect 27 108 715 109
rect 27 106 134 108
rect 136 106 388 108
rect 390 106 715 108
rect 27 103 715 106
rect 24 102 69 103
rect 24 100 25 102
rect 27 101 69 102
rect 71 102 715 103
rect 71 101 106 102
rect 27 100 106 101
rect 108 100 177 102
rect 179 100 242 102
rect 244 100 295 102
rect 297 101 363 102
rect 297 100 330 101
rect 24 99 330 100
rect 332 100 363 101
rect 365 100 409 102
rect 411 100 454 102
rect 456 101 712 102
rect 456 100 527 101
rect 332 99 527 100
rect 529 99 592 101
rect 594 100 712 101
rect 714 100 715 102
rect 594 99 715 100
rect 27 96 715 99
rect 27 94 44 96
rect 46 94 387 96
rect 389 94 715 96
rect 27 93 715 94
rect 31 87 43 88
rect 31 85 33 87
rect 35 85 43 87
rect 31 82 43 85
rect 31 80 35 82
rect 31 78 33 80
rect 31 55 35 78
rect 143 83 156 87
rect 244 83 257 87
rect 374 87 386 88
rect 345 83 358 87
rect 55 78 77 80
rect 151 81 156 83
rect 151 79 152 81
rect 154 79 156 81
rect 55 76 74 78
rect 76 76 77 78
rect 55 74 67 76
rect 31 53 36 55
rect 31 51 33 53
rect 35 51 36 53
rect 31 46 36 51
rect 47 64 51 72
rect 47 62 59 64
rect 47 60 50 62
rect 52 61 59 62
rect 52 60 55 61
rect 47 59 55 60
rect 57 59 59 61
rect 47 58 59 59
rect 63 62 67 74
rect 65 60 67 62
rect 63 58 67 60
rect 71 71 77 76
rect 71 69 74 71
rect 76 69 77 71
rect 71 67 77 69
rect 31 44 33 46
rect 35 44 36 46
rect 31 42 36 44
rect 71 47 75 67
rect 87 70 125 71
rect 87 68 88 70
rect 90 68 125 70
rect 87 67 125 68
rect 120 64 125 67
rect 95 62 110 63
rect 95 60 99 62
rect 101 60 106 62
rect 108 60 110 62
rect 95 59 110 60
rect 120 62 128 64
rect 120 60 125 62
rect 127 60 128 62
rect 104 50 108 59
rect 120 58 128 60
rect 151 74 156 79
rect 151 72 152 74
rect 154 72 156 74
rect 151 70 156 72
rect 71 46 93 47
rect 71 44 74 46
rect 76 44 93 46
rect 71 43 93 44
rect 152 48 156 70
rect 151 46 156 48
rect 151 44 152 46
rect 154 44 156 46
rect 151 42 156 44
rect 172 78 178 80
rect 252 81 257 83
rect 252 79 253 81
rect 255 79 257 81
rect 172 76 175 78
rect 177 76 178 78
rect 172 71 178 76
rect 172 69 175 71
rect 177 69 178 71
rect 172 67 178 69
rect 172 53 176 67
rect 188 70 226 71
rect 188 68 189 70
rect 191 68 226 70
rect 188 67 226 68
rect 221 64 226 67
rect 196 62 211 63
rect 196 60 200 62
rect 202 60 207 62
rect 209 60 211 62
rect 196 59 211 60
rect 221 62 229 64
rect 221 60 226 62
rect 228 60 229 62
rect 172 51 173 53
rect 175 51 176 53
rect 172 47 176 51
rect 205 53 209 59
rect 221 58 229 60
rect 252 74 257 79
rect 252 72 253 74
rect 255 72 257 74
rect 252 70 257 72
rect 253 61 257 70
rect 253 59 254 61
rect 256 59 257 61
rect 205 51 206 53
rect 208 51 209 53
rect 205 50 209 51
rect 172 46 194 47
rect 172 44 175 46
rect 177 44 194 46
rect 172 43 194 44
rect 253 48 257 59
rect 252 46 257 48
rect 252 44 253 46
rect 255 44 257 46
rect 252 42 257 44
rect 273 78 279 80
rect 353 81 358 83
rect 353 79 354 81
rect 356 79 358 81
rect 273 76 276 78
rect 278 76 279 78
rect 273 71 279 76
rect 273 69 276 71
rect 278 69 279 71
rect 273 67 279 69
rect 273 53 277 67
rect 289 70 327 71
rect 289 68 290 70
rect 292 68 327 70
rect 289 67 327 68
rect 322 64 327 67
rect 297 62 312 63
rect 297 60 301 62
rect 303 60 308 62
rect 310 60 312 62
rect 297 59 312 60
rect 322 62 330 64
rect 322 60 327 62
rect 329 60 330 62
rect 306 58 310 59
rect 322 58 330 60
rect 273 51 274 53
rect 276 51 277 53
rect 306 56 307 58
rect 309 56 310 58
rect 273 47 277 51
rect 306 50 310 56
rect 353 74 358 79
rect 353 72 354 74
rect 356 72 358 74
rect 353 70 358 72
rect 273 46 295 47
rect 273 44 276 46
rect 278 44 295 46
rect 273 43 295 44
rect 354 48 358 70
rect 353 46 358 48
rect 353 44 354 46
rect 356 44 358 46
rect 353 42 358 44
rect 374 85 376 87
rect 378 85 386 87
rect 374 82 386 85
rect 374 80 378 82
rect 374 78 376 80
rect 374 58 378 78
rect 498 83 511 87
rect 599 83 612 87
rect 698 83 711 87
rect 374 56 375 58
rect 377 56 378 58
rect 374 55 378 56
rect 398 78 432 80
rect 506 81 511 83
rect 506 79 507 81
rect 509 79 511 81
rect 398 76 429 78
rect 431 76 432 78
rect 398 74 410 76
rect 374 53 379 55
rect 374 51 376 53
rect 378 51 379 53
rect 374 46 379 51
rect 390 64 394 72
rect 390 62 402 64
rect 390 60 393 62
rect 395 61 402 62
rect 395 60 398 61
rect 390 59 398 60
rect 400 59 402 61
rect 390 58 402 59
rect 406 62 410 74
rect 408 60 410 62
rect 406 58 410 60
rect 426 71 432 76
rect 426 69 429 71
rect 431 69 432 71
rect 426 67 432 69
rect 374 44 376 46
rect 378 44 379 46
rect 374 42 379 44
rect 426 47 430 67
rect 442 70 480 71
rect 442 68 443 70
rect 445 68 480 70
rect 442 67 480 68
rect 475 64 480 67
rect 450 62 465 63
rect 450 60 454 62
rect 456 60 461 62
rect 463 60 465 62
rect 450 59 465 60
rect 475 62 483 64
rect 475 60 480 62
rect 482 60 483 62
rect 459 50 463 59
rect 475 58 483 60
rect 506 74 511 79
rect 506 72 507 74
rect 509 72 511 74
rect 506 70 511 72
rect 426 46 448 47
rect 426 44 429 46
rect 431 44 448 46
rect 426 43 448 44
rect 507 48 511 70
rect 506 46 511 48
rect 506 44 507 46
rect 509 44 511 46
rect 506 42 511 44
rect 527 78 533 80
rect 607 81 612 83
rect 607 79 608 81
rect 610 79 612 81
rect 527 76 530 78
rect 532 76 533 78
rect 527 71 533 76
rect 527 69 530 71
rect 532 69 533 71
rect 527 67 533 69
rect 527 53 531 67
rect 543 70 581 71
rect 543 68 544 70
rect 546 68 581 70
rect 543 67 581 68
rect 576 64 581 67
rect 551 62 566 63
rect 551 60 555 62
rect 557 60 562 62
rect 564 60 566 62
rect 551 59 566 60
rect 576 62 584 64
rect 576 60 581 62
rect 583 60 584 62
rect 527 51 528 53
rect 530 51 531 53
rect 527 47 531 51
rect 560 53 564 59
rect 576 58 584 60
rect 607 74 612 79
rect 607 72 608 74
rect 610 72 612 74
rect 607 70 612 72
rect 608 61 612 70
rect 608 59 609 61
rect 611 59 612 61
rect 560 51 561 53
rect 563 51 564 53
rect 560 50 564 51
rect 527 46 549 47
rect 527 44 530 46
rect 532 44 549 46
rect 527 43 549 44
rect 608 48 612 59
rect 607 46 612 48
rect 607 44 608 46
rect 610 44 612 46
rect 607 42 612 44
rect 626 78 632 80
rect 706 81 711 83
rect 706 79 707 81
rect 709 79 711 81
rect 626 76 629 78
rect 631 76 632 78
rect 626 71 632 76
rect 626 69 629 71
rect 631 69 632 71
rect 626 67 632 69
rect 626 53 630 67
rect 642 70 680 71
rect 642 68 643 70
rect 645 68 680 70
rect 642 67 680 68
rect 675 64 680 67
rect 650 62 665 63
rect 650 60 651 62
rect 653 60 654 62
rect 656 60 661 62
rect 663 60 665 62
rect 650 59 665 60
rect 675 62 683 64
rect 675 60 680 62
rect 682 60 683 62
rect 626 51 627 53
rect 629 51 630 53
rect 626 47 630 51
rect 659 50 663 59
rect 675 58 683 60
rect 706 74 711 79
rect 706 72 707 74
rect 709 72 711 74
rect 706 70 711 72
rect 626 46 648 47
rect 626 44 629 46
rect 631 44 648 46
rect 626 43 648 44
rect 707 48 711 70
rect 706 46 711 48
rect 706 44 707 46
rect 709 44 711 46
rect 706 42 711 44
rect 27 36 715 37
rect 27 34 60 36
rect 62 34 403 36
rect 405 34 715 36
rect 27 32 28 34
rect 30 32 89 34
rect 91 32 153 34
rect 155 32 217 34
rect 219 32 280 34
rect 282 32 316 34
rect 318 32 347 34
rect 349 32 388 34
rect 390 32 419 34
rect 421 32 476 34
rect 478 32 566 34
rect 568 32 669 34
rect 671 32 712 34
rect 714 32 715 34
rect 27 29 715 32
<< alu2 >>
rect 362 390 366 391
rect 362 388 363 390
rect 365 388 366 390
rect 67 387 71 388
rect 362 387 366 388
rect 408 390 412 391
rect 408 388 409 390
rect 411 388 412 390
rect 408 387 412 388
rect 453 390 457 391
rect 453 388 454 390
rect 456 388 457 390
rect 453 387 457 388
rect 526 390 530 391
rect 526 388 527 390
rect 529 388 530 390
rect 526 387 530 388
rect 712 387 716 388
rect 27 386 31 387
rect 27 384 28 386
rect 30 384 31 386
rect 67 385 68 387
rect 70 385 71 387
rect 67 384 71 385
rect 105 386 109 387
rect 105 384 106 386
rect 108 384 109 386
rect 27 383 31 384
rect 105 383 109 384
rect 176 386 180 387
rect 176 384 177 386
rect 179 384 180 386
rect 176 383 180 384
rect 241 386 245 387
rect 241 384 242 386
rect 244 384 245 386
rect 241 383 245 384
rect 294 386 298 387
rect 294 384 295 386
rect 297 384 298 386
rect 294 383 298 384
rect 329 386 333 387
rect 329 384 330 386
rect 332 384 333 386
rect 329 383 333 384
rect 591 386 595 387
rect 591 384 592 386
rect 594 384 595 386
rect 712 385 713 387
rect 715 385 716 387
rect 712 384 716 385
rect 591 383 595 384
rect 360 382 560 383
rect 360 380 361 382
rect 363 380 557 382
rect 559 380 560 382
rect 360 379 560 380
rect 62 374 131 375
rect 62 372 63 374
rect 65 372 128 374
rect 130 372 131 374
rect 62 371 131 372
rect 273 374 342 375
rect 273 372 274 374
rect 276 372 339 374
rect 341 372 342 374
rect 273 371 342 372
rect 443 374 512 375
rect 443 372 444 374
rect 446 372 509 374
rect 511 372 512 374
rect 443 371 512 372
rect 578 374 647 375
rect 578 372 579 374
rect 581 372 644 374
rect 646 372 647 374
rect 578 371 647 372
rect 71 366 503 367
rect 71 364 72 366
rect 74 364 500 366
rect 502 364 503 366
rect 71 363 503 364
rect 40 358 75 359
rect 40 356 41 358
rect 43 356 72 358
rect 74 356 75 358
rect 40 355 75 356
rect 127 358 131 359
rect 127 356 128 358
rect 130 356 131 358
rect 127 355 131 356
rect 273 358 277 359
rect 273 356 274 358
rect 276 356 277 358
rect 273 355 277 356
rect 329 358 364 359
rect 329 356 330 358
rect 332 356 361 358
rect 363 356 364 358
rect 329 355 364 356
rect 443 358 447 359
rect 443 356 444 358
rect 446 356 447 358
rect 443 355 447 356
rect 499 358 534 359
rect 499 356 500 358
rect 502 356 531 358
rect 533 356 534 358
rect 499 355 534 356
rect 556 358 591 359
rect 556 356 557 358
rect 559 356 588 358
rect 590 356 591 358
rect 556 355 591 356
rect 643 358 647 359
rect 643 356 644 358
rect 646 356 647 358
rect 643 355 647 356
rect 38 350 366 351
rect 38 348 39 350
rect 41 348 363 350
rect 365 348 366 350
rect 38 347 366 348
rect 492 349 598 350
rect 492 347 493 349
rect 495 347 595 349
rect 597 347 598 349
rect 492 346 598 347
rect 38 341 42 342
rect 38 339 39 341
rect 41 339 42 341
rect 38 338 42 339
rect 78 341 82 342
rect 78 339 79 341
rect 81 339 82 341
rect 78 338 82 339
rect 144 341 148 342
rect 144 339 145 341
rect 147 339 148 341
rect 144 338 148 339
rect 256 341 260 342
rect 256 339 257 341
rect 259 339 260 341
rect 256 338 260 339
rect 322 341 326 342
rect 322 339 323 341
rect 325 339 326 341
rect 322 338 326 339
rect 362 341 366 342
rect 362 339 363 341
rect 365 339 366 341
rect 362 338 366 339
rect 426 341 430 342
rect 426 339 427 341
rect 429 339 430 341
rect 426 338 430 339
rect 492 341 496 342
rect 492 339 493 341
rect 495 339 496 341
rect 492 338 496 339
rect 532 341 536 342
rect 532 339 533 341
rect 535 339 536 341
rect 532 338 536 339
rect 554 341 558 342
rect 554 339 555 341
rect 557 339 558 341
rect 554 338 558 339
rect 594 341 598 342
rect 594 339 595 341
rect 597 339 598 341
rect 594 338 598 339
rect 660 341 664 342
rect 660 339 661 341
rect 663 339 664 341
rect 660 338 664 339
rect 129 334 133 335
rect 102 333 110 334
rect 102 331 103 333
rect 105 331 107 333
rect 109 331 110 333
rect 129 332 130 334
rect 132 332 133 334
rect 129 331 133 332
rect 191 334 200 335
rect 191 332 192 334
rect 194 332 197 334
rect 199 332 200 334
rect 191 331 200 332
rect 209 334 213 335
rect 209 332 210 334
rect 212 332 213 334
rect 209 331 213 332
rect 271 334 275 335
rect 379 334 383 335
rect 271 332 272 334
rect 274 332 275 334
rect 271 331 275 332
rect 294 333 302 334
rect 294 331 295 333
rect 297 331 299 333
rect 301 331 302 333
rect 379 332 380 334
rect 382 332 383 334
rect 379 331 383 332
rect 441 334 445 335
rect 645 334 649 335
rect 441 332 442 334
rect 444 332 445 334
rect 441 331 445 332
rect 464 333 472 334
rect 464 331 465 333
rect 467 331 469 333
rect 471 331 472 333
rect 102 330 110 331
rect 294 330 302 331
rect 464 330 472 331
rect 618 333 626 334
rect 618 331 619 333
rect 621 331 623 333
rect 625 331 626 333
rect 645 332 646 334
rect 648 332 649 334
rect 645 331 649 332
rect 618 330 626 331
rect 27 318 31 319
rect 27 316 28 318
rect 30 316 31 318
rect 27 315 31 316
rect 88 318 92 319
rect 88 316 89 318
rect 91 316 92 318
rect 88 315 92 316
rect 152 318 156 319
rect 152 316 153 318
rect 155 316 156 318
rect 152 315 156 316
rect 216 318 220 319
rect 216 316 217 318
rect 219 316 220 318
rect 216 315 220 316
rect 279 318 283 319
rect 279 316 280 318
rect 282 316 283 318
rect 279 315 283 316
rect 314 318 318 319
rect 314 316 315 318
rect 317 316 318 318
rect 314 315 318 316
rect 346 318 350 319
rect 346 316 347 318
rect 349 316 350 318
rect 346 315 350 316
rect 387 318 391 319
rect 387 316 388 318
rect 390 316 391 318
rect 387 315 391 316
rect 418 318 422 319
rect 418 316 419 318
rect 421 316 422 318
rect 418 315 422 316
rect 475 318 479 319
rect 475 316 476 318
rect 478 316 479 318
rect 475 315 479 316
rect 565 318 569 319
rect 565 316 566 318
rect 568 316 569 318
rect 565 315 569 316
rect 668 318 672 319
rect 668 316 669 318
rect 671 316 672 318
rect 668 315 672 316
rect 712 318 716 319
rect 712 316 713 318
rect 715 316 716 318
rect 712 315 716 316
rect 102 303 148 304
rect 102 301 103 303
rect 105 301 145 303
rect 147 301 148 303
rect 102 300 148 301
rect 256 303 302 304
rect 256 301 257 303
rect 259 301 299 303
rect 301 301 302 303
rect 256 300 302 301
rect 426 303 472 304
rect 426 301 427 303
rect 429 301 469 303
rect 471 301 472 303
rect 426 300 472 301
rect 618 303 664 304
rect 618 301 619 303
rect 621 301 661 303
rect 663 301 664 303
rect 618 300 664 301
rect 38 295 42 296
rect 38 293 39 295
rect 41 293 42 295
rect 38 292 42 293
rect 78 295 326 296
rect 78 293 79 295
rect 81 293 323 295
rect 325 293 326 295
rect 78 292 326 293
rect 362 295 366 296
rect 492 295 496 296
rect 362 293 363 295
rect 365 293 366 295
rect 362 292 366 293
rect 418 294 463 295
rect 418 292 419 294
rect 421 292 460 294
rect 462 292 463 294
rect 492 293 493 295
rect 495 293 496 295
rect 492 292 496 293
rect 532 295 558 296
rect 532 293 533 295
rect 535 293 555 295
rect 557 293 558 295
rect 532 292 558 293
rect 594 295 598 296
rect 594 293 595 295
rect 597 293 598 295
rect 594 292 598 293
rect 418 291 463 292
rect 59 286 67 287
rect 59 284 60 286
rect 62 284 64 286
rect 66 284 67 286
rect 59 283 67 284
rect 129 286 139 287
rect 129 284 130 286
rect 132 284 136 286
rect 138 284 139 286
rect 129 283 139 284
rect 208 286 261 287
rect 208 284 209 286
rect 211 284 258 286
rect 260 284 261 286
rect 208 283 261 284
rect 265 286 275 287
rect 265 284 266 286
rect 268 284 272 286
rect 274 284 275 286
rect 265 283 275 284
rect 435 286 445 287
rect 435 284 436 286
rect 438 284 442 286
rect 444 284 445 286
rect 435 283 445 284
rect 507 286 522 287
rect 507 284 508 286
rect 510 284 519 286
rect 521 284 522 286
rect 507 283 522 284
rect 645 286 655 287
rect 645 284 646 286
rect 648 284 652 286
rect 654 284 655 286
rect 645 283 655 284
rect 40 278 75 279
rect 40 276 41 278
rect 43 276 68 278
rect 70 276 72 278
rect 74 276 75 278
rect 40 275 75 276
rect 106 278 131 279
rect 106 276 107 278
rect 109 276 128 278
rect 130 276 131 278
rect 106 275 131 276
rect 168 278 222 279
rect 168 276 169 278
rect 171 276 219 278
rect 221 276 222 278
rect 168 275 222 276
rect 273 278 298 279
rect 273 276 274 278
rect 276 276 295 278
rect 297 276 298 278
rect 273 275 298 276
rect 329 278 364 279
rect 329 276 330 278
rect 332 276 361 278
rect 363 276 364 278
rect 329 275 364 276
rect 443 278 468 279
rect 443 276 444 278
rect 446 276 465 278
rect 467 276 468 278
rect 443 275 468 276
rect 499 278 534 279
rect 499 276 500 278
rect 502 276 531 278
rect 533 276 534 278
rect 499 275 534 276
rect 556 278 591 279
rect 556 276 557 278
rect 559 276 588 278
rect 590 276 591 278
rect 556 275 591 276
rect 622 278 647 279
rect 622 276 623 278
rect 625 276 644 278
rect 646 276 647 278
rect 622 275 647 276
rect 369 274 383 275
rect 369 272 370 274
rect 372 272 380 274
rect 382 272 383 274
rect 369 271 383 272
rect 113 270 117 271
rect 113 268 114 270
rect 116 268 117 270
rect 218 270 291 271
rect 218 268 219 270
rect 221 268 288 270
rect 290 268 291 270
rect 113 267 117 268
rect 187 267 195 268
rect 187 265 188 267
rect 190 265 192 267
rect 194 265 195 267
rect 187 264 195 265
rect 209 267 213 268
rect 218 267 291 268
rect 613 270 633 271
rect 613 268 614 270
rect 616 268 630 270
rect 632 268 633 270
rect 613 267 633 268
rect 209 265 210 267
rect 212 265 213 267
rect 209 264 213 265
rect 338 265 342 266
rect 338 263 339 265
rect 341 263 342 265
rect 338 262 342 263
rect 360 265 560 266
rect 360 263 361 265
rect 363 263 557 265
rect 559 263 560 265
rect 360 262 560 263
rect 699 262 703 263
rect 699 260 700 262
rect 702 260 703 262
rect 699 259 703 260
rect 67 257 503 258
rect 67 255 68 257
rect 70 255 500 257
rect 502 255 503 257
rect 67 254 503 255
rect 712 247 716 248
rect 67 246 71 247
rect 27 245 31 246
rect 27 243 28 245
rect 30 243 31 245
rect 67 244 68 246
rect 70 244 71 246
rect 67 243 71 244
rect 105 246 109 247
rect 105 244 106 246
rect 108 244 109 246
rect 105 243 109 244
rect 176 246 180 247
rect 176 244 177 246
rect 179 244 180 246
rect 176 243 180 244
rect 241 246 245 247
rect 241 244 242 246
rect 244 244 245 246
rect 241 243 245 244
rect 294 246 298 247
rect 408 246 412 247
rect 294 244 295 246
rect 297 244 298 246
rect 294 243 298 244
rect 329 245 333 246
rect 329 243 330 245
rect 332 243 333 245
rect 27 242 31 243
rect 329 242 333 243
rect 361 245 365 246
rect 361 243 362 245
rect 364 243 365 245
rect 408 244 409 246
rect 411 244 412 246
rect 408 243 412 244
rect 453 246 457 247
rect 453 244 454 246
rect 456 244 457 246
rect 453 243 457 244
rect 526 245 530 246
rect 526 243 527 245
rect 529 243 530 245
rect 361 242 365 243
rect 526 242 530 243
rect 591 245 595 246
rect 591 243 592 245
rect 594 243 595 245
rect 712 245 713 247
rect 715 245 716 247
rect 712 244 716 245
rect 591 242 595 243
rect 152 230 294 231
rect 152 228 153 230
rect 155 228 291 230
rect 293 228 294 230
rect 152 227 294 228
rect 338 230 647 231
rect 338 228 339 230
rect 341 228 644 230
rect 646 228 647 230
rect 338 227 647 228
rect 257 222 447 223
rect 257 220 258 222
rect 260 220 444 222
rect 446 220 447 222
rect 257 219 447 220
rect 518 222 655 223
rect 518 220 519 222
rect 521 220 652 222
rect 654 220 655 222
rect 518 219 655 220
rect 121 214 164 215
rect 121 212 122 214
rect 124 212 161 214
rect 163 212 164 214
rect 121 211 164 212
rect 209 214 213 215
rect 209 212 210 214
rect 212 212 213 214
rect 209 211 213 212
rect 290 214 294 215
rect 290 212 291 214
rect 293 212 294 214
rect 290 211 294 212
rect 318 214 422 215
rect 318 212 319 214
rect 321 212 419 214
rect 421 212 422 214
rect 318 211 422 212
rect 443 214 447 215
rect 443 212 444 214
rect 446 212 447 214
rect 443 211 447 212
rect 544 214 548 215
rect 544 212 545 214
rect 547 212 548 214
rect 544 211 548 212
rect 643 214 647 215
rect 643 212 644 214
rect 646 212 647 214
rect 643 211 647 212
rect 206 206 379 207
rect 461 206 465 207
rect 651 206 655 207
rect 52 205 56 206
rect 52 203 53 205
rect 55 203 56 205
rect 52 202 56 203
rect 113 205 125 206
rect 113 203 114 205
rect 116 203 122 205
rect 124 203 125 205
rect 206 204 207 206
rect 209 204 376 206
rect 378 204 379 206
rect 206 203 379 204
rect 398 205 402 206
rect 398 203 399 205
rect 401 203 402 205
rect 113 202 125 203
rect 160 198 268 199
rect 398 198 402 203
rect 461 204 462 206
rect 464 205 613 206
rect 464 204 610 205
rect 461 203 610 204
rect 612 203 613 205
rect 651 204 652 206
rect 654 204 655 206
rect 651 203 655 204
rect 461 202 613 203
rect 104 197 116 198
rect 104 195 105 197
rect 107 195 113 197
rect 115 195 116 197
rect 160 196 161 198
rect 163 196 265 198
rect 267 196 268 198
rect 160 195 268 196
rect 307 197 311 198
rect 307 195 308 197
rect 310 195 311 197
rect 104 194 116 195
rect 307 194 311 195
rect 398 197 532 198
rect 398 195 529 197
rect 531 195 532 197
rect 398 194 532 195
rect 561 197 631 198
rect 561 195 562 197
rect 564 195 628 197
rect 630 195 631 197
rect 561 194 631 195
rect 32 190 36 191
rect 32 188 33 190
rect 35 188 36 190
rect 32 187 36 188
rect 144 190 178 191
rect 144 188 145 190
rect 147 188 175 190
rect 177 188 178 190
rect 144 187 178 188
rect 205 190 256 191
rect 354 190 358 191
rect 660 190 711 191
rect 205 188 207 190
rect 209 188 253 190
rect 255 188 256 190
rect 205 187 256 188
rect 264 189 322 190
rect 264 187 265 189
rect 267 187 319 189
rect 321 187 322 189
rect 354 188 355 190
rect 357 188 358 190
rect 354 187 358 188
rect 504 189 508 190
rect 504 187 505 189
rect 507 187 508 189
rect 660 188 661 190
rect 663 188 708 190
rect 710 188 711 190
rect 660 187 711 188
rect 264 186 322 187
rect 504 186 508 187
rect 379 181 548 182
rect 379 179 380 181
rect 382 179 545 181
rect 547 179 548 181
rect 379 178 548 179
rect 24 174 28 175
rect 152 174 156 175
rect 24 172 25 174
rect 27 172 28 174
rect 24 171 28 172
rect 88 173 92 174
rect 88 171 89 173
rect 91 171 92 173
rect 152 172 153 174
rect 155 172 156 174
rect 152 171 156 172
rect 216 174 220 175
rect 216 172 217 174
rect 219 172 220 174
rect 216 171 220 172
rect 279 174 283 175
rect 279 172 280 174
rect 282 172 283 174
rect 279 171 283 172
rect 315 174 319 175
rect 315 172 316 174
rect 318 172 319 174
rect 315 171 319 172
rect 346 174 350 175
rect 565 174 569 175
rect 346 172 347 174
rect 349 172 350 174
rect 346 171 350 172
rect 387 173 391 174
rect 387 171 388 173
rect 390 171 391 173
rect 88 170 92 171
rect 387 170 391 171
rect 418 173 422 174
rect 418 171 419 173
rect 421 171 422 173
rect 418 170 422 171
rect 475 173 479 174
rect 475 171 476 173
rect 478 171 479 173
rect 565 172 566 174
rect 568 172 569 174
rect 565 171 569 172
rect 668 174 672 175
rect 668 172 669 174
rect 671 172 672 174
rect 668 171 672 172
rect 712 174 716 175
rect 712 172 713 174
rect 715 172 716 174
rect 712 171 716 172
rect 475 170 479 171
rect 50 158 54 159
rect 50 156 51 158
rect 53 156 54 158
rect 50 155 54 156
rect 112 158 116 159
rect 112 156 113 158
rect 115 156 116 158
rect 112 155 116 156
rect 307 158 341 159
rect 307 156 308 158
rect 310 156 338 158
rect 340 156 341 158
rect 307 155 341 156
rect 122 151 126 152
rect 65 150 123 151
rect 65 148 66 150
rect 68 149 123 150
rect 125 149 126 151
rect 68 148 126 149
rect 206 151 210 152
rect 398 151 532 152
rect 206 149 207 151
rect 209 149 210 151
rect 206 148 210 149
rect 254 150 326 151
rect 254 148 255 150
rect 257 148 323 150
rect 325 148 326 150
rect 65 147 126 148
rect 254 147 326 148
rect 398 149 529 151
rect 531 149 532 151
rect 398 148 532 149
rect 561 151 631 152
rect 561 149 562 151
rect 564 149 628 151
rect 630 149 631 151
rect 561 148 631 149
rect 660 151 664 152
rect 660 149 661 151
rect 663 149 664 151
rect 660 148 664 149
rect 144 143 148 144
rect 398 143 402 148
rect 144 141 145 143
rect 147 141 148 143
rect 144 140 148 141
rect 226 142 373 143
rect 226 140 227 142
rect 229 140 370 142
rect 372 140 373 142
rect 398 141 399 143
rect 401 141 402 143
rect 398 140 402 141
rect 461 143 613 144
rect 461 142 610 143
rect 461 140 462 142
rect 464 141 610 142
rect 612 141 613 143
rect 464 140 613 141
rect 226 139 373 140
rect 461 139 465 140
rect 578 135 617 136
rect 82 134 172 135
rect 82 132 83 134
rect 85 132 169 134
rect 171 132 172 134
rect 82 131 172 132
rect 339 134 379 135
rect 339 132 340 134
rect 342 132 376 134
rect 378 132 379 134
rect 339 131 379 132
rect 477 134 508 135
rect 477 132 478 134
rect 480 132 505 134
rect 507 132 508 134
rect 578 133 579 135
rect 581 133 614 135
rect 616 133 617 135
rect 578 132 617 133
rect 677 134 703 135
rect 677 132 678 134
rect 680 132 700 134
rect 702 132 703 134
rect 477 131 508 132
rect 677 131 703 132
rect 283 118 287 119
rect 283 116 284 118
rect 286 116 287 118
rect 283 115 287 116
rect 283 110 654 111
rect 283 108 284 110
rect 286 108 651 110
rect 653 108 654 110
rect 283 107 654 108
rect 68 103 72 104
rect 24 102 28 103
rect 24 100 25 102
rect 27 100 28 102
rect 68 101 69 103
rect 71 101 72 103
rect 68 100 72 101
rect 105 102 109 103
rect 105 100 106 102
rect 108 100 109 102
rect 24 99 28 100
rect 105 99 109 100
rect 176 102 180 103
rect 176 100 177 102
rect 179 100 180 102
rect 176 99 180 100
rect 241 102 245 103
rect 241 100 242 102
rect 244 100 245 102
rect 241 99 245 100
rect 294 102 298 103
rect 362 102 366 103
rect 294 100 295 102
rect 297 100 298 102
rect 294 99 298 100
rect 329 101 333 102
rect 329 99 330 101
rect 332 99 333 101
rect 362 100 363 102
rect 365 100 366 102
rect 362 99 366 100
rect 408 102 412 103
rect 408 100 409 102
rect 411 100 412 102
rect 408 99 412 100
rect 453 102 457 103
rect 711 102 715 103
rect 453 100 454 102
rect 456 100 457 102
rect 453 99 457 100
rect 526 101 530 102
rect 526 99 527 101
rect 529 99 530 101
rect 329 98 333 99
rect 526 98 530 99
rect 591 101 595 102
rect 591 99 592 101
rect 594 99 595 101
rect 711 100 712 102
rect 714 100 715 102
rect 711 99 715 100
rect 591 98 595 99
rect 354 92 446 93
rect 354 90 355 92
rect 357 90 443 92
rect 445 90 446 92
rect 354 89 446 90
rect 60 86 350 87
rect 60 84 61 86
rect 63 85 350 86
rect 63 84 646 85
rect 60 83 643 84
rect 346 82 643 83
rect 645 82 646 84
rect 346 81 646 82
rect 187 78 293 79
rect 187 76 188 78
rect 190 76 290 78
rect 292 76 293 78
rect 187 75 293 76
rect 32 70 91 71
rect 32 68 33 70
rect 35 68 88 70
rect 90 68 91 70
rect 32 67 91 68
rect 121 70 192 71
rect 121 68 122 70
rect 124 68 189 70
rect 191 68 192 70
rect 121 67 192 68
rect 289 70 293 71
rect 289 68 290 70
rect 292 68 293 70
rect 289 67 293 68
rect 442 70 446 71
rect 442 68 443 70
rect 445 68 446 70
rect 442 67 446 68
rect 543 70 547 71
rect 543 68 544 70
rect 546 68 547 70
rect 543 67 547 68
rect 642 70 646 71
rect 642 68 643 70
rect 645 68 646 70
rect 642 67 646 68
rect 105 62 109 63
rect 460 62 464 63
rect 650 62 654 63
rect 54 61 58 62
rect 54 59 55 61
rect 57 59 58 61
rect 54 54 58 59
rect 105 60 106 62
rect 108 61 257 62
rect 108 60 254 61
rect 105 59 254 60
rect 256 59 257 61
rect 397 61 401 62
rect 397 59 398 61
rect 400 59 401 61
rect 105 58 257 59
rect 306 58 378 59
rect 306 56 307 58
rect 309 56 375 58
rect 377 56 378 58
rect 306 55 378 56
rect 397 54 401 59
rect 460 60 461 62
rect 463 61 612 62
rect 463 60 609 61
rect 460 59 609 60
rect 611 59 612 61
rect 650 60 651 62
rect 653 60 654 62
rect 650 59 654 60
rect 460 58 612 59
rect 54 53 176 54
rect 54 51 173 53
rect 175 51 176 53
rect 54 50 176 51
rect 205 53 277 54
rect 205 51 206 53
rect 208 51 274 53
rect 276 51 277 53
rect 205 50 277 51
rect 397 53 531 54
rect 397 51 528 53
rect 530 51 531 53
rect 397 50 531 51
rect 560 53 630 54
rect 560 51 561 53
rect 563 51 627 53
rect 629 51 630 53
rect 560 50 630 51
rect 196 45 547 46
rect 196 43 197 45
rect 199 43 544 45
rect 546 43 547 45
rect 196 42 547 43
rect 27 34 31 35
rect 27 32 28 34
rect 30 32 31 34
rect 27 31 31 32
rect 88 34 92 35
rect 88 32 89 34
rect 91 32 92 34
rect 88 31 92 32
rect 152 34 156 35
rect 152 32 153 34
rect 155 32 156 34
rect 152 31 156 32
rect 216 34 220 35
rect 216 32 217 34
rect 219 32 220 34
rect 216 31 220 32
rect 279 34 283 35
rect 279 32 280 34
rect 282 32 283 34
rect 279 31 283 32
rect 315 34 319 35
rect 315 32 316 34
rect 318 32 319 34
rect 315 31 319 32
rect 346 34 350 35
rect 346 32 347 34
rect 349 32 350 34
rect 346 31 350 32
rect 387 34 391 35
rect 387 32 388 34
rect 390 32 391 34
rect 387 31 391 32
rect 418 34 422 35
rect 418 32 419 34
rect 421 32 422 34
rect 418 31 422 32
rect 475 34 479 35
rect 475 32 476 34
rect 478 32 479 34
rect 475 31 479 32
rect 565 34 569 35
rect 565 32 566 34
rect 568 32 569 34
rect 565 31 569 32
rect 668 34 672 35
rect 668 32 669 34
rect 671 32 672 34
rect 668 31 672 32
rect 711 34 715 35
rect 711 32 712 34
rect 714 32 715 34
rect 711 31 715 32
<< alu3 >>
rect 362 390 366 391
rect 362 388 363 390
rect 365 388 366 390
rect 67 387 71 388
rect 362 387 366 388
rect 408 390 412 391
rect 408 388 409 390
rect 411 388 412 390
rect 408 387 412 388
rect 453 390 457 391
rect 453 388 454 390
rect 456 388 457 390
rect 453 387 457 388
rect 526 390 530 391
rect 526 388 527 390
rect 529 388 530 390
rect 526 387 530 388
rect 712 387 716 388
rect 27 386 31 387
rect 27 384 28 386
rect 30 384 31 386
rect 67 385 68 387
rect 70 385 71 387
rect 67 384 71 385
rect 105 386 109 387
rect 105 384 106 386
rect 108 384 109 386
rect 27 383 31 384
rect 105 383 109 384
rect 176 386 180 387
rect 176 384 177 386
rect 179 384 180 386
rect 176 383 180 384
rect 241 386 245 387
rect 241 384 242 386
rect 244 384 245 386
rect 241 383 245 384
rect 294 386 298 387
rect 294 384 295 386
rect 297 384 298 386
rect 294 383 298 384
rect 329 386 333 387
rect 329 384 330 386
rect 332 384 333 386
rect 329 383 333 384
rect 591 386 595 387
rect 591 384 592 386
rect 594 384 595 386
rect 712 385 713 387
rect 715 385 716 387
rect 712 384 716 385
rect 591 383 595 384
rect 360 382 364 383
rect 360 380 361 382
rect 363 380 364 382
rect 127 374 131 375
rect 127 372 128 374
rect 130 372 131 374
rect 71 366 75 367
rect 71 364 72 366
rect 74 364 75 366
rect 71 358 75 364
rect 71 356 72 358
rect 74 356 75 358
rect 71 355 75 356
rect 127 358 131 372
rect 127 356 128 358
rect 130 356 131 358
rect 127 355 131 356
rect 273 374 277 375
rect 273 372 274 374
rect 276 372 277 374
rect 273 358 277 372
rect 273 356 274 358
rect 276 356 277 358
rect 273 355 277 356
rect 360 358 364 380
rect 556 382 560 383
rect 556 380 557 382
rect 559 380 560 382
rect 360 356 361 358
rect 363 356 364 358
rect 360 355 364 356
rect 443 374 447 375
rect 443 372 444 374
rect 446 372 447 374
rect 443 358 447 372
rect 443 356 444 358
rect 446 356 447 358
rect 443 355 447 356
rect 499 366 503 367
rect 499 364 500 366
rect 502 364 503 366
rect 499 358 503 364
rect 499 356 500 358
rect 502 356 503 358
rect 499 355 503 356
rect 556 358 560 380
rect 556 356 557 358
rect 559 356 560 358
rect 556 355 560 356
rect 643 374 647 375
rect 643 372 644 374
rect 646 372 647 374
rect 643 358 647 372
rect 643 356 644 358
rect 646 356 647 358
rect 643 355 647 356
rect 38 350 42 351
rect 38 348 39 350
rect 41 348 42 350
rect 38 341 42 348
rect 362 350 366 351
rect 362 348 363 350
rect 365 348 366 350
rect 38 339 39 341
rect 41 339 42 341
rect 27 318 31 319
rect 27 316 28 318
rect 30 316 31 318
rect 27 315 31 316
rect 38 295 42 339
rect 38 293 39 295
rect 41 293 42 295
rect 38 292 42 293
rect 78 341 82 342
rect 78 339 79 341
rect 81 339 82 341
rect 78 295 82 339
rect 144 341 148 342
rect 144 339 145 341
rect 147 339 148 341
rect 129 334 133 335
rect 106 333 110 334
rect 106 331 107 333
rect 109 331 110 333
rect 88 318 92 319
rect 88 316 89 318
rect 91 316 92 318
rect 88 315 92 316
rect 78 293 79 295
rect 81 293 82 295
rect 78 292 82 293
rect 59 286 63 287
rect 59 284 60 286
rect 62 284 63 286
rect 27 245 31 246
rect 27 243 28 245
rect 30 243 31 245
rect 27 242 31 243
rect 59 214 63 284
rect 67 278 71 279
rect 67 276 68 278
rect 70 276 71 278
rect 67 257 71 276
rect 106 278 110 331
rect 129 332 130 334
rect 132 332 133 334
rect 129 286 133 332
rect 144 303 148 339
rect 256 341 260 342
rect 256 339 257 341
rect 259 339 260 341
rect 196 334 200 335
rect 196 332 197 334
rect 199 332 200 334
rect 152 318 156 319
rect 152 316 153 318
rect 155 316 156 318
rect 152 315 156 316
rect 144 301 145 303
rect 147 301 148 303
rect 144 300 148 301
rect 129 284 130 286
rect 132 284 133 286
rect 129 283 133 284
rect 106 276 107 278
rect 109 276 110 278
rect 106 275 110 276
rect 168 278 172 279
rect 168 276 169 278
rect 171 276 172 278
rect 67 255 68 257
rect 70 255 71 257
rect 67 254 71 255
rect 113 270 117 271
rect 113 268 114 270
rect 116 268 117 270
rect 67 246 71 247
rect 67 244 68 246
rect 70 244 71 246
rect 67 243 71 244
rect 105 246 109 247
rect 105 244 106 246
rect 108 244 109 246
rect 105 243 109 244
rect 59 210 64 214
rect 50 205 56 206
rect 50 203 53 205
rect 55 203 56 205
rect 50 202 56 203
rect 32 190 36 191
rect 32 188 33 190
rect 35 188 36 190
rect 24 174 28 175
rect 24 172 25 174
rect 27 172 28 174
rect 24 171 28 172
rect 24 102 28 103
rect 24 100 25 102
rect 27 100 28 102
rect 24 99 28 100
rect 32 70 36 188
rect 50 158 54 202
rect 50 156 51 158
rect 53 156 54 158
rect 50 155 54 156
rect 60 86 64 210
rect 113 205 117 268
rect 160 214 164 215
rect 160 212 161 214
rect 163 212 164 214
rect 113 203 114 205
rect 116 203 117 205
rect 113 202 117 203
rect 121 205 125 206
rect 121 203 122 205
rect 124 203 125 205
rect 112 197 116 198
rect 112 195 113 197
rect 115 195 116 197
rect 88 173 92 174
rect 88 171 89 173
rect 91 171 92 173
rect 88 170 92 171
rect 112 158 116 195
rect 112 156 113 158
rect 115 156 116 158
rect 112 155 116 156
rect 68 103 72 104
rect 68 101 69 103
rect 71 101 72 103
rect 68 100 72 101
rect 105 102 109 103
rect 105 100 106 102
rect 108 100 109 102
rect 105 99 109 100
rect 60 84 61 86
rect 63 84 64 86
rect 60 83 64 84
rect 32 68 33 70
rect 35 68 36 70
rect 32 67 36 68
rect 121 70 125 203
rect 160 198 164 212
rect 160 196 161 198
rect 163 196 164 198
rect 160 195 164 196
rect 144 190 148 191
rect 144 188 145 190
rect 147 188 148 190
rect 144 143 148 188
rect 152 174 156 175
rect 152 172 153 174
rect 155 172 156 174
rect 152 171 156 172
rect 144 141 145 143
rect 147 141 148 143
rect 144 140 148 141
rect 168 134 172 276
rect 187 267 191 268
rect 187 265 188 267
rect 190 265 191 267
rect 176 246 180 247
rect 176 244 177 246
rect 179 244 180 246
rect 176 243 180 244
rect 168 132 169 134
rect 171 132 172 134
rect 168 131 172 132
rect 176 102 180 103
rect 176 100 177 102
rect 179 100 180 102
rect 176 99 180 100
rect 187 78 191 265
rect 187 76 188 78
rect 190 76 191 78
rect 187 75 191 76
rect 121 68 122 70
rect 124 68 125 70
rect 121 67 125 68
rect 196 45 200 332
rect 208 334 213 335
rect 208 332 210 334
rect 212 332 213 334
rect 208 331 213 332
rect 208 286 212 331
rect 216 318 220 319
rect 216 316 217 318
rect 219 316 220 318
rect 216 315 220 316
rect 256 303 260 339
rect 322 341 326 342
rect 322 339 323 341
rect 325 339 326 341
rect 256 301 257 303
rect 259 301 260 303
rect 256 300 260 301
rect 271 334 275 335
rect 271 332 272 334
rect 274 332 275 334
rect 208 284 209 286
rect 211 284 212 286
rect 208 283 212 284
rect 257 286 261 287
rect 257 284 258 286
rect 260 284 261 286
rect 218 278 222 279
rect 218 276 219 278
rect 221 276 222 278
rect 218 270 222 276
rect 218 268 219 270
rect 221 268 222 270
rect 209 267 213 268
rect 218 267 222 268
rect 209 265 210 267
rect 212 265 213 267
rect 209 214 213 265
rect 241 246 245 247
rect 241 244 242 246
rect 244 244 245 246
rect 241 243 245 244
rect 257 222 261 284
rect 271 286 275 332
rect 294 333 298 334
rect 294 331 295 333
rect 297 331 298 333
rect 279 318 283 319
rect 279 316 280 318
rect 282 316 283 318
rect 279 315 283 316
rect 271 284 272 286
rect 274 284 275 286
rect 271 283 275 284
rect 294 278 298 331
rect 314 318 318 319
rect 314 316 315 318
rect 317 316 318 318
rect 314 315 318 316
rect 322 295 326 339
rect 362 341 366 348
rect 492 349 496 350
rect 492 347 493 349
rect 495 347 496 349
rect 362 339 363 341
rect 365 339 366 341
rect 346 318 350 319
rect 346 316 347 318
rect 349 316 350 318
rect 346 315 350 316
rect 322 293 323 295
rect 325 293 326 295
rect 322 292 326 293
rect 362 295 366 339
rect 426 341 430 342
rect 426 339 427 341
rect 429 339 430 341
rect 362 293 363 295
rect 365 293 366 295
rect 362 292 366 293
rect 379 334 383 335
rect 379 332 380 334
rect 382 332 383 334
rect 294 276 295 278
rect 297 276 298 278
rect 294 275 298 276
rect 360 278 364 279
rect 360 276 361 278
rect 363 276 364 278
rect 338 265 342 266
rect 338 263 339 265
rect 341 263 342 265
rect 294 246 298 247
rect 294 244 295 246
rect 297 244 298 246
rect 294 243 298 244
rect 329 245 333 246
rect 329 243 330 245
rect 332 243 333 245
rect 329 242 333 243
rect 257 220 258 222
rect 260 220 261 222
rect 257 219 261 220
rect 290 230 294 231
rect 290 228 291 230
rect 293 228 294 230
rect 209 212 210 214
rect 212 212 213 214
rect 209 211 213 212
rect 290 214 294 228
rect 338 230 342 263
rect 360 265 364 276
rect 360 263 361 265
rect 363 263 364 265
rect 360 262 364 263
rect 369 274 373 275
rect 369 272 370 274
rect 372 272 373 274
rect 361 245 365 246
rect 361 243 362 245
rect 364 243 365 245
rect 361 242 365 243
rect 338 228 339 230
rect 341 228 342 230
rect 338 227 342 228
rect 290 212 291 214
rect 293 212 294 214
rect 290 211 294 212
rect 318 214 322 215
rect 318 212 319 214
rect 321 212 322 214
rect 264 198 268 199
rect 264 196 265 198
rect 267 196 268 198
rect 206 190 210 191
rect 206 188 207 190
rect 209 188 210 190
rect 206 151 210 188
rect 264 189 268 196
rect 264 187 265 189
rect 267 187 268 189
rect 264 186 268 187
rect 307 197 311 198
rect 307 195 308 197
rect 310 195 311 197
rect 216 174 220 175
rect 216 172 217 174
rect 219 172 220 174
rect 216 171 220 172
rect 279 174 283 175
rect 279 172 280 174
rect 282 172 283 174
rect 279 171 283 172
rect 307 158 311 195
rect 318 189 322 212
rect 318 187 319 189
rect 321 187 322 189
rect 318 186 322 187
rect 354 190 358 191
rect 354 188 355 190
rect 357 188 358 190
rect 315 174 319 175
rect 315 172 316 174
rect 318 172 319 174
rect 315 171 319 172
rect 346 174 350 175
rect 346 172 347 174
rect 349 172 350 174
rect 346 171 350 172
rect 307 156 308 158
rect 310 156 311 158
rect 307 155 311 156
rect 206 149 207 151
rect 209 149 210 151
rect 206 148 210 149
rect 283 118 287 119
rect 283 116 284 118
rect 286 116 287 118
rect 283 110 287 116
rect 283 108 284 110
rect 286 108 287 110
rect 283 107 287 108
rect 241 102 245 103
rect 241 100 242 102
rect 244 100 245 102
rect 241 99 245 100
rect 294 102 298 103
rect 294 100 295 102
rect 297 100 298 102
rect 294 99 298 100
rect 329 101 333 102
rect 329 99 330 101
rect 332 99 333 101
rect 329 98 333 99
rect 354 92 358 188
rect 369 142 373 272
rect 379 181 383 332
rect 387 318 391 319
rect 387 316 388 318
rect 390 316 391 318
rect 387 315 391 316
rect 418 318 422 319
rect 418 316 419 318
rect 421 316 422 318
rect 418 315 422 316
rect 426 303 430 339
rect 492 341 496 347
rect 594 349 598 350
rect 594 347 595 349
rect 597 347 598 349
rect 492 339 493 341
rect 495 339 496 341
rect 426 301 427 303
rect 429 301 430 303
rect 426 300 430 301
rect 441 334 445 335
rect 441 332 442 334
rect 444 332 445 334
rect 418 294 422 295
rect 418 292 419 294
rect 421 292 422 294
rect 408 246 412 247
rect 408 244 409 246
rect 411 244 412 246
rect 408 243 412 244
rect 418 214 422 292
rect 441 286 445 332
rect 441 284 442 286
rect 444 284 445 286
rect 441 283 445 284
rect 464 333 468 334
rect 464 331 465 333
rect 467 331 468 333
rect 464 278 468 331
rect 475 318 479 319
rect 475 316 476 318
rect 478 316 479 318
rect 475 315 479 316
rect 492 295 496 339
rect 492 293 493 295
rect 495 293 496 295
rect 492 292 496 293
rect 532 341 536 342
rect 532 339 533 341
rect 535 339 536 341
rect 532 295 536 339
rect 532 293 533 295
rect 535 293 536 295
rect 532 292 536 293
rect 554 341 558 342
rect 554 339 555 341
rect 557 339 558 341
rect 554 295 558 339
rect 594 341 598 347
rect 594 339 595 341
rect 597 339 598 341
rect 565 318 569 319
rect 565 316 566 318
rect 568 316 569 318
rect 565 315 569 316
rect 554 293 555 295
rect 557 293 558 295
rect 554 292 558 293
rect 594 295 598 339
rect 660 341 664 342
rect 660 339 661 341
rect 663 339 664 341
rect 645 334 649 335
rect 594 293 595 295
rect 597 293 598 295
rect 594 292 598 293
rect 622 333 626 334
rect 622 331 623 333
rect 625 331 626 333
rect 518 286 522 287
rect 518 284 519 286
rect 521 284 522 286
rect 464 276 465 278
rect 467 276 468 278
rect 464 275 468 276
rect 499 278 503 279
rect 499 276 500 278
rect 502 276 503 278
rect 499 257 503 276
rect 499 255 500 257
rect 502 255 503 257
rect 499 254 503 255
rect 453 246 457 247
rect 453 244 454 246
rect 456 244 457 246
rect 453 243 457 244
rect 418 212 419 214
rect 421 212 422 214
rect 418 211 422 212
rect 443 222 447 223
rect 443 220 444 222
rect 446 220 447 222
rect 443 214 447 220
rect 518 222 522 284
rect 556 278 560 279
rect 556 276 557 278
rect 559 276 560 278
rect 556 265 560 276
rect 622 278 626 331
rect 645 332 646 334
rect 648 332 649 334
rect 645 286 649 332
rect 660 303 664 339
rect 668 318 672 319
rect 668 316 669 318
rect 671 316 672 318
rect 668 315 672 316
rect 712 318 716 319
rect 712 316 713 318
rect 715 316 716 318
rect 712 315 716 316
rect 660 301 661 303
rect 663 301 664 303
rect 660 300 664 301
rect 645 284 646 286
rect 648 284 649 286
rect 645 283 649 284
rect 622 276 623 278
rect 625 276 626 278
rect 622 275 626 276
rect 556 263 557 265
rect 559 263 560 265
rect 556 262 560 263
rect 613 270 617 271
rect 613 268 614 270
rect 616 268 617 270
rect 526 245 530 246
rect 526 243 527 245
rect 529 243 530 245
rect 526 242 530 243
rect 591 245 595 246
rect 591 243 592 245
rect 594 243 595 245
rect 591 242 595 243
rect 518 220 519 222
rect 521 220 522 222
rect 518 219 522 220
rect 443 212 444 214
rect 446 212 447 214
rect 443 211 447 212
rect 544 214 548 215
rect 544 212 545 214
rect 547 212 548 214
rect 379 179 380 181
rect 382 179 383 181
rect 379 178 383 179
rect 504 189 508 190
rect 504 187 505 189
rect 507 187 508 189
rect 387 173 391 174
rect 387 171 388 173
rect 390 171 391 173
rect 387 170 391 171
rect 418 173 422 174
rect 418 171 419 173
rect 421 171 422 173
rect 418 170 422 171
rect 475 173 479 174
rect 475 171 476 173
rect 478 171 479 173
rect 475 170 479 171
rect 369 140 370 142
rect 372 140 373 142
rect 369 139 373 140
rect 504 134 508 187
rect 544 181 548 212
rect 544 179 545 181
rect 547 179 548 181
rect 544 178 548 179
rect 565 174 569 175
rect 565 172 566 174
rect 568 172 569 174
rect 565 171 569 172
rect 504 132 505 134
rect 507 132 508 134
rect 613 135 617 268
rect 699 262 703 263
rect 699 260 700 262
rect 702 260 703 262
rect 643 230 647 231
rect 643 228 644 230
rect 646 228 647 230
rect 643 214 647 228
rect 643 212 644 214
rect 646 212 647 214
rect 643 211 647 212
rect 651 222 655 223
rect 651 220 652 222
rect 654 220 655 222
rect 651 206 655 220
rect 651 204 652 206
rect 654 204 655 206
rect 651 203 655 204
rect 660 190 664 191
rect 660 188 661 190
rect 663 188 664 190
rect 660 151 664 188
rect 668 174 672 175
rect 668 172 669 174
rect 671 172 672 174
rect 668 171 672 172
rect 660 149 661 151
rect 663 149 664 151
rect 660 148 664 149
rect 613 133 614 135
rect 616 133 617 135
rect 613 132 617 133
rect 699 134 703 260
rect 712 247 716 248
rect 712 245 713 247
rect 715 245 716 247
rect 712 244 716 245
rect 712 174 716 175
rect 712 172 713 174
rect 715 172 716 174
rect 712 171 716 172
rect 699 132 700 134
rect 702 132 703 134
rect 504 131 508 132
rect 699 131 703 132
rect 650 110 654 111
rect 650 108 651 110
rect 653 108 654 110
rect 362 102 366 103
rect 362 100 363 102
rect 365 100 366 102
rect 362 99 366 100
rect 408 102 412 103
rect 408 100 409 102
rect 411 100 412 102
rect 408 99 412 100
rect 453 102 457 103
rect 453 100 454 102
rect 456 100 457 102
rect 453 99 457 100
rect 526 101 530 102
rect 526 99 527 101
rect 529 99 530 101
rect 526 98 530 99
rect 591 101 595 102
rect 591 99 592 101
rect 594 99 595 101
rect 591 98 595 99
rect 354 90 355 92
rect 357 90 358 92
rect 354 89 358 90
rect 442 92 446 93
rect 442 90 443 92
rect 445 90 446 92
rect 289 78 293 79
rect 289 76 290 78
rect 292 76 293 78
rect 289 70 293 76
rect 289 68 290 70
rect 292 68 293 70
rect 289 67 293 68
rect 442 70 446 90
rect 642 84 646 85
rect 642 82 643 84
rect 645 82 646 84
rect 442 68 443 70
rect 445 68 446 70
rect 442 67 446 68
rect 543 70 547 71
rect 543 68 544 70
rect 546 68 547 70
rect 196 43 197 45
rect 199 43 200 45
rect 196 42 200 43
rect 543 45 547 68
rect 642 70 646 82
rect 642 68 643 70
rect 645 68 646 70
rect 642 67 646 68
rect 650 62 654 108
rect 711 102 715 103
rect 711 100 712 102
rect 714 100 715 102
rect 711 99 715 100
rect 650 60 651 62
rect 653 60 654 62
rect 650 59 654 60
rect 543 43 544 45
rect 546 43 547 45
rect 543 42 547 43
rect 27 34 31 35
rect 27 32 28 34
rect 30 32 31 34
rect 27 31 31 32
rect 88 34 92 35
rect 88 32 89 34
rect 91 32 92 34
rect 88 31 92 32
rect 152 34 156 35
rect 152 32 153 34
rect 155 32 156 34
rect 152 31 156 32
rect 216 34 220 35
rect 216 32 217 34
rect 219 32 220 34
rect 216 31 220 32
rect 279 34 283 35
rect 279 32 280 34
rect 282 32 283 34
rect 279 31 283 32
rect 315 34 319 35
rect 315 32 316 34
rect 318 32 319 34
rect 315 31 319 32
rect 346 34 350 35
rect 346 32 347 34
rect 349 32 350 34
rect 346 31 350 32
rect 387 34 391 35
rect 387 32 388 34
rect 390 32 391 34
rect 387 31 391 32
rect 418 34 422 35
rect 418 32 419 34
rect 421 32 422 34
rect 418 31 422 32
rect 475 34 479 35
rect 475 32 476 34
rect 478 32 479 34
rect 475 31 479 32
rect 565 34 569 35
rect 565 32 566 34
rect 568 32 569 34
rect 565 31 569 32
rect 668 34 672 35
rect 668 32 669 34
rect 671 32 672 34
rect 668 31 672 32
rect 711 34 715 35
rect 711 32 712 34
rect 714 32 715 34
rect 711 31 715 32
<< alu4 >>
rect 0 413 8 414
rect 0 411 5 413
rect 7 411 8 413
rect 0 318 8 411
rect 88 413 92 414
rect 88 411 89 413
rect 91 411 92 413
rect 0 316 5 318
rect 7 316 8 318
rect 0 174 8 316
rect 0 172 5 174
rect 7 172 8 174
rect 0 34 8 172
rect 0 32 5 34
rect 7 32 8 34
rect 0 7 8 32
rect 12 401 20 402
rect 12 399 17 401
rect 19 399 20 401
rect 12 386 20 399
rect 67 401 71 402
rect 67 399 68 401
rect 70 399 71 401
rect 67 387 71 399
rect 12 384 17 386
rect 19 384 20 386
rect 12 245 20 384
rect 27 386 31 387
rect 27 384 28 386
rect 30 384 31 386
rect 27 383 31 384
rect 67 385 68 387
rect 70 385 71 387
rect 27 318 31 319
rect 27 316 28 318
rect 30 316 31 318
rect 27 315 31 316
rect 67 246 71 385
rect 12 243 17 245
rect 19 243 20 245
rect 12 102 20 243
rect 27 245 31 246
rect 27 243 28 245
rect 30 243 31 245
rect 27 242 31 243
rect 67 244 68 246
rect 70 244 71 246
rect 24 174 28 175
rect 24 172 25 174
rect 27 172 28 174
rect 24 171 28 172
rect 67 104 71 244
rect 88 318 92 411
rect 152 413 156 414
rect 152 411 153 413
rect 155 411 156 413
rect 88 316 89 318
rect 91 316 92 318
rect 88 173 92 316
rect 88 171 89 173
rect 91 171 92 173
rect 67 103 72 104
rect 12 100 17 102
rect 19 100 20 102
rect 12 19 20 100
rect 24 102 28 103
rect 24 100 25 102
rect 27 100 28 102
rect 24 99 28 100
rect 67 101 69 103
rect 71 101 72 103
rect 67 100 72 101
rect 27 34 31 35
rect 27 32 28 34
rect 30 32 31 34
rect 27 31 31 32
rect 12 17 17 19
rect 19 17 20 19
rect 12 16 20 17
rect 67 19 71 100
rect 67 17 68 19
rect 70 17 71 19
rect 67 16 71 17
rect 88 34 92 171
rect 88 32 89 34
rect 91 32 92 34
rect 0 5 5 7
rect 7 5 8 7
rect 0 4 8 5
rect 88 7 92 32
rect 105 401 109 402
rect 105 399 106 401
rect 108 399 109 401
rect 105 386 109 399
rect 105 384 106 386
rect 108 384 109 386
rect 105 246 109 384
rect 105 244 106 246
rect 108 244 109 246
rect 105 102 109 244
rect 105 100 106 102
rect 108 100 109 102
rect 105 19 109 100
rect 105 17 106 19
rect 108 17 109 19
rect 105 16 109 17
rect 152 318 156 411
rect 216 413 220 414
rect 216 411 217 413
rect 219 411 220 413
rect 152 316 153 318
rect 155 316 156 318
rect 152 174 156 316
rect 152 172 153 174
rect 155 172 156 174
rect 152 34 156 172
rect 152 32 153 34
rect 155 32 156 34
rect 88 5 89 7
rect 91 5 92 7
rect 88 4 92 5
rect 152 7 156 32
rect 176 401 180 402
rect 176 399 177 401
rect 179 399 180 401
rect 176 386 180 399
rect 176 384 177 386
rect 179 384 180 386
rect 176 246 180 384
rect 176 244 177 246
rect 179 244 180 246
rect 176 102 180 244
rect 176 100 177 102
rect 179 100 180 102
rect 176 19 180 100
rect 176 17 177 19
rect 179 17 180 19
rect 176 16 180 17
rect 216 318 220 411
rect 279 413 283 414
rect 279 411 280 413
rect 282 411 283 413
rect 216 316 217 318
rect 219 316 220 318
rect 216 174 220 316
rect 216 172 217 174
rect 219 172 220 174
rect 216 34 220 172
rect 216 32 217 34
rect 219 32 220 34
rect 152 5 153 7
rect 155 5 156 7
rect 152 4 156 5
rect 216 7 220 32
rect 241 401 245 402
rect 241 399 242 401
rect 244 399 245 401
rect 241 386 245 399
rect 241 384 242 386
rect 244 384 245 386
rect 241 246 245 384
rect 241 244 242 246
rect 244 244 245 246
rect 241 102 245 244
rect 241 100 242 102
rect 244 100 245 102
rect 241 19 245 100
rect 241 17 242 19
rect 244 17 245 19
rect 241 16 245 17
rect 279 318 283 411
rect 315 413 319 414
rect 315 411 316 413
rect 318 411 319 413
rect 279 316 280 318
rect 282 316 283 318
rect 279 174 283 316
rect 279 172 280 174
rect 282 172 283 174
rect 279 34 283 172
rect 279 32 280 34
rect 282 32 283 34
rect 216 5 217 7
rect 219 5 220 7
rect 216 4 220 5
rect 279 7 283 32
rect 294 401 298 402
rect 294 399 295 401
rect 297 399 298 401
rect 294 386 298 399
rect 294 384 295 386
rect 297 384 298 386
rect 294 246 298 384
rect 315 319 319 411
rect 346 413 350 414
rect 346 411 347 413
rect 349 411 350 413
rect 314 318 319 319
rect 314 316 315 318
rect 317 316 319 318
rect 314 315 319 316
rect 294 244 295 246
rect 297 244 298 246
rect 294 102 298 244
rect 294 100 295 102
rect 297 100 298 102
rect 294 19 298 100
rect 294 17 295 19
rect 297 17 298 19
rect 294 16 298 17
rect 315 174 319 315
rect 315 172 316 174
rect 318 172 319 174
rect 315 34 319 172
rect 315 32 316 34
rect 318 32 319 34
rect 279 5 280 7
rect 282 5 283 7
rect 279 4 283 5
rect 315 7 319 32
rect 329 401 333 402
rect 329 399 330 401
rect 332 399 333 401
rect 329 386 333 399
rect 329 384 330 386
rect 332 384 333 386
rect 329 245 333 384
rect 329 243 330 245
rect 332 243 333 245
rect 329 101 333 243
rect 329 99 330 101
rect 332 99 333 101
rect 329 19 333 99
rect 329 17 330 19
rect 332 17 333 19
rect 329 16 333 17
rect 346 318 350 411
rect 387 413 391 414
rect 387 411 388 413
rect 390 411 391 413
rect 346 316 347 318
rect 349 316 350 318
rect 346 174 350 316
rect 362 401 366 402
rect 362 399 363 401
rect 365 399 366 401
rect 362 390 366 399
rect 362 388 363 390
rect 365 388 366 390
rect 362 246 366 388
rect 361 245 366 246
rect 361 243 362 245
rect 364 243 366 245
rect 361 242 366 243
rect 346 172 347 174
rect 349 172 350 174
rect 346 34 350 172
rect 346 32 347 34
rect 349 32 350 34
rect 315 5 316 7
rect 318 5 319 7
rect 315 4 319 5
rect 346 7 350 32
rect 362 102 366 242
rect 362 100 363 102
rect 365 100 366 102
rect 362 19 366 100
rect 362 17 363 19
rect 365 17 366 19
rect 362 16 366 17
rect 387 318 391 411
rect 418 413 422 414
rect 418 411 419 413
rect 421 411 422 413
rect 387 316 388 318
rect 390 316 391 318
rect 387 173 391 316
rect 387 171 388 173
rect 390 171 391 173
rect 387 34 391 171
rect 387 32 388 34
rect 390 32 391 34
rect 346 5 347 7
rect 349 5 350 7
rect 346 4 350 5
rect 387 7 391 32
rect 408 401 412 402
rect 408 399 409 401
rect 411 399 412 401
rect 408 390 412 399
rect 408 388 409 390
rect 411 388 412 390
rect 408 246 412 388
rect 408 244 409 246
rect 411 244 412 246
rect 408 102 412 244
rect 408 100 409 102
rect 411 100 412 102
rect 408 19 412 100
rect 408 17 409 19
rect 411 17 412 19
rect 408 16 412 17
rect 418 318 422 411
rect 475 413 479 414
rect 475 411 476 413
rect 478 411 479 413
rect 418 316 419 318
rect 421 316 422 318
rect 418 173 422 316
rect 418 171 419 173
rect 421 171 422 173
rect 418 34 422 171
rect 418 32 419 34
rect 421 32 422 34
rect 387 5 388 7
rect 390 5 391 7
rect 387 4 391 5
rect 418 7 422 32
rect 453 401 457 402
rect 453 399 454 401
rect 456 399 457 401
rect 453 390 457 399
rect 453 388 454 390
rect 456 388 457 390
rect 453 246 457 388
rect 453 244 454 246
rect 456 244 457 246
rect 453 102 457 244
rect 453 100 454 102
rect 456 100 457 102
rect 453 19 457 100
rect 453 17 454 19
rect 456 17 457 19
rect 453 16 457 17
rect 475 318 479 411
rect 565 413 569 414
rect 565 411 566 413
rect 568 411 569 413
rect 475 316 476 318
rect 478 316 479 318
rect 475 173 479 316
rect 475 171 476 173
rect 478 171 479 173
rect 475 34 479 171
rect 475 32 476 34
rect 478 32 479 34
rect 418 5 419 7
rect 421 5 422 7
rect 418 4 422 5
rect 475 7 479 32
rect 526 401 530 402
rect 526 399 527 401
rect 529 399 530 401
rect 526 390 530 399
rect 526 388 527 390
rect 529 388 530 390
rect 526 245 530 388
rect 526 243 527 245
rect 529 243 530 245
rect 526 101 530 243
rect 526 99 527 101
rect 529 99 530 101
rect 526 19 530 99
rect 526 17 527 19
rect 529 17 530 19
rect 526 16 530 17
rect 565 318 569 411
rect 668 413 672 414
rect 668 411 669 413
rect 671 411 672 413
rect 565 316 566 318
rect 568 316 569 318
rect 565 174 569 316
rect 565 172 566 174
rect 568 172 569 174
rect 565 34 569 172
rect 565 32 566 34
rect 568 32 569 34
rect 475 5 476 7
rect 478 5 479 7
rect 475 4 479 5
rect 565 7 569 32
rect 591 401 595 402
rect 591 399 592 401
rect 594 399 595 401
rect 591 386 595 399
rect 591 384 592 386
rect 594 384 595 386
rect 591 245 595 384
rect 591 243 592 245
rect 594 243 595 245
rect 591 101 595 243
rect 591 99 592 101
rect 594 99 595 101
rect 591 19 595 99
rect 591 17 592 19
rect 594 17 595 19
rect 591 16 595 17
rect 668 318 672 411
rect 734 413 742 414
rect 734 411 735 413
rect 737 411 742 413
rect 722 401 730 402
rect 722 399 723 401
rect 725 399 730 401
rect 712 387 716 388
rect 712 385 713 387
rect 715 385 716 387
rect 712 384 716 385
rect 722 387 730 399
rect 722 385 723 387
rect 725 385 730 387
rect 668 316 669 318
rect 671 316 672 318
rect 668 174 672 316
rect 712 318 716 319
rect 712 316 713 318
rect 715 316 716 318
rect 712 315 716 316
rect 712 247 716 248
rect 712 245 713 247
rect 715 245 716 247
rect 712 244 716 245
rect 722 247 730 385
rect 722 245 723 247
rect 725 245 730 247
rect 668 172 669 174
rect 671 172 672 174
rect 668 34 672 172
rect 712 174 716 175
rect 712 172 713 174
rect 715 172 716 174
rect 712 171 716 172
rect 711 102 715 103
rect 711 100 712 102
rect 714 100 715 102
rect 711 99 715 100
rect 722 102 730 245
rect 722 100 723 102
rect 725 100 730 102
rect 668 32 669 34
rect 671 32 672 34
rect 565 5 566 7
rect 568 5 569 7
rect 565 4 569 5
rect 668 7 672 32
rect 711 34 715 35
rect 711 32 712 34
rect 714 32 715 34
rect 711 31 715 32
rect 722 19 730 100
rect 722 17 723 19
rect 725 17 730 19
rect 722 16 730 17
rect 734 318 742 411
rect 734 316 735 318
rect 737 316 742 318
rect 734 174 742 316
rect 734 172 735 174
rect 737 172 742 174
rect 734 34 742 172
rect 734 32 735 34
rect 737 32 742 34
rect 668 5 669 7
rect 671 5 672 7
rect 668 4 672 5
rect 734 7 742 32
rect 734 5 735 7
rect 737 5 742 7
rect 734 4 742 5
<< alu5 >>
rect 4 413 738 418
rect 4 411 5 413
rect 7 411 89 413
rect 91 411 153 413
rect 155 411 217 413
rect 219 411 280 413
rect 282 411 316 413
rect 318 411 347 413
rect 349 411 388 413
rect 390 411 419 413
rect 421 411 476 413
rect 478 411 566 413
rect 568 411 669 413
rect 671 411 735 413
rect 737 411 738 413
rect 4 410 738 411
rect 16 401 726 406
rect 16 399 17 401
rect 19 399 68 401
rect 70 399 106 401
rect 108 399 177 401
rect 179 399 242 401
rect 244 399 295 401
rect 297 399 330 401
rect 332 399 363 401
rect 365 399 409 401
rect 411 399 454 401
rect 456 399 527 401
rect 529 399 592 401
rect 594 399 723 401
rect 725 399 726 401
rect 16 398 726 399
rect 712 387 726 388
rect 16 386 31 387
rect 16 384 17 386
rect 19 384 28 386
rect 30 384 31 386
rect 712 385 713 387
rect 715 385 723 387
rect 725 385 726 387
rect 712 384 726 385
rect 16 383 31 384
rect 4 318 31 319
rect 4 316 5 318
rect 7 316 28 318
rect 30 316 31 318
rect 4 315 31 316
rect 712 318 738 319
rect 712 316 713 318
rect 715 316 735 318
rect 737 316 738 318
rect 712 315 738 316
rect 712 247 726 248
rect 16 245 31 246
rect 16 243 17 245
rect 19 243 28 245
rect 30 243 31 245
rect 712 245 713 247
rect 715 245 723 247
rect 725 245 726 247
rect 712 244 726 245
rect 16 242 31 243
rect 4 174 28 175
rect 4 172 5 174
rect 7 172 25 174
rect 27 172 28 174
rect 4 171 28 172
rect 712 174 738 175
rect 712 172 713 174
rect 715 172 735 174
rect 737 172 738 174
rect 712 171 738 172
rect 16 102 28 103
rect 16 100 17 102
rect 19 100 25 102
rect 27 100 28 102
rect 16 99 28 100
rect 711 102 726 103
rect 711 100 712 102
rect 714 100 723 102
rect 725 100 726 102
rect 711 99 726 100
rect 4 34 31 35
rect 4 32 5 34
rect 7 32 28 34
rect 30 32 31 34
rect 4 31 31 32
rect 711 34 738 35
rect 711 32 712 34
rect 714 32 735 34
rect 737 32 738 34
rect 711 31 738 32
rect 16 19 726 20
rect 16 17 17 19
rect 19 17 68 19
rect 70 17 106 19
rect 108 17 177 19
rect 179 17 242 19
rect 244 17 295 19
rect 297 17 330 19
rect 332 17 363 19
rect 365 17 409 19
rect 411 17 454 19
rect 456 17 527 19
rect 529 17 592 19
rect 594 17 723 19
rect 725 17 726 19
rect 16 12 726 17
rect 4 7 738 8
rect 4 5 5 7
rect 7 5 89 7
rect 91 5 153 7
rect 155 5 217 7
rect 219 5 280 7
rect 282 5 316 7
rect 318 5 347 7
rect 349 5 388 7
rect 390 5 419 7
rect 421 5 476 7
rect 478 5 566 7
rect 568 5 669 7
rect 671 5 735 7
rect 737 5 738 7
rect 4 0 738 5
<< ptie >>
rect 56 176 66 182
rect 400 180 410 182
rect 400 178 404 180
rect 406 178 410 180
rect 400 176 410 178
rect 146 168 156 170
rect 146 166 150 168
rect 152 166 156 168
rect 146 164 156 166
rect 400 168 410 170
rect 400 166 404 168
rect 406 166 410 168
rect 400 164 410 166
rect 56 36 66 38
rect 56 34 60 36
rect 62 34 66 36
rect 56 32 66 34
rect 399 36 409 38
rect 399 34 403 36
rect 405 34 409 36
rect 399 32 409 34
<< nmos >>
rect 38 330 40 343
rect 45 330 47 343
rect 58 329 60 343
rect 78 330 80 343
rect 85 330 87 343
rect 98 329 100 343
rect 119 323 121 337
rect 130 323 132 343
rect 137 323 139 343
rect 157 329 159 343
rect 167 329 169 343
rect 177 326 179 336
rect 187 323 189 336
rect 215 323 217 336
rect 225 326 227 336
rect 235 329 237 343
rect 245 329 247 343
rect 265 323 267 343
rect 272 323 274 343
rect 283 323 285 337
rect 304 329 306 343
rect 317 330 319 343
rect 324 330 326 343
rect 344 329 346 343
rect 357 330 359 343
rect 364 330 366 343
rect 385 323 387 336
rect 395 326 397 336
rect 405 329 407 343
rect 415 329 417 343
rect 435 323 437 343
rect 442 323 444 343
rect 453 323 455 337
rect 474 329 476 343
rect 487 330 489 343
rect 494 330 496 343
rect 514 329 516 343
rect 527 330 529 343
rect 534 330 536 343
rect 554 330 556 343
rect 561 330 563 343
rect 574 329 576 343
rect 594 330 596 343
rect 601 330 603 343
rect 614 329 616 343
rect 635 323 637 337
rect 646 323 648 343
rect 653 323 655 343
rect 673 329 675 343
rect 683 329 685 343
rect 693 326 695 336
rect 703 323 705 336
rect 38 291 40 304
rect 45 291 47 304
rect 58 291 60 305
rect 78 291 80 304
rect 85 291 87 304
rect 98 291 100 305
rect 119 297 121 311
rect 130 291 132 311
rect 137 291 139 311
rect 157 291 159 305
rect 167 291 169 305
rect 177 298 179 308
rect 187 298 189 311
rect 215 298 217 311
rect 225 298 227 308
rect 235 291 237 305
rect 245 291 247 305
rect 265 291 267 311
rect 272 291 274 311
rect 283 297 285 311
rect 304 291 306 305
rect 317 291 319 304
rect 324 291 326 304
rect 344 291 346 305
rect 357 291 359 304
rect 364 291 366 304
rect 385 298 387 311
rect 395 298 397 308
rect 405 291 407 305
rect 415 291 417 305
rect 435 291 437 311
rect 442 291 444 311
rect 453 297 455 311
rect 474 291 476 305
rect 487 291 489 304
rect 494 291 496 304
rect 514 291 516 305
rect 527 291 529 304
rect 534 291 536 304
rect 554 291 556 304
rect 561 291 563 304
rect 574 291 576 305
rect 594 291 596 304
rect 601 291 603 304
rect 614 291 616 305
rect 635 297 637 311
rect 646 291 648 311
rect 653 291 655 311
rect 673 291 675 305
rect 683 291 685 305
rect 693 298 695 308
rect 703 298 705 311
rect 38 185 40 199
rect 48 186 50 194
rect 58 188 60 196
rect 79 179 81 193
rect 90 179 92 199
rect 97 179 99 199
rect 117 185 119 199
rect 127 185 129 199
rect 137 182 139 192
rect 147 179 149 192
rect 180 179 182 193
rect 191 179 193 199
rect 198 179 200 199
rect 218 185 220 199
rect 228 185 230 199
rect 238 182 240 192
rect 248 179 250 192
rect 282 179 284 193
rect 293 179 295 199
rect 300 179 302 199
rect 320 185 322 199
rect 330 185 332 199
rect 340 182 342 192
rect 350 179 352 192
rect 382 185 384 199
rect 392 186 394 194
rect 402 188 404 196
rect 435 179 437 193
rect 446 179 448 199
rect 453 179 455 199
rect 473 185 475 199
rect 483 185 485 199
rect 493 182 495 192
rect 503 179 505 192
rect 536 179 538 193
rect 547 179 549 199
rect 554 179 556 199
rect 574 185 576 199
rect 584 185 586 199
rect 594 182 596 192
rect 604 179 606 192
rect 635 179 637 193
rect 646 179 648 199
rect 653 179 655 199
rect 673 185 675 199
rect 683 185 685 199
rect 693 182 695 192
rect 703 179 705 192
rect 40 153 42 167
rect 51 147 53 167
rect 58 147 60 167
rect 78 147 80 161
rect 88 147 90 161
rect 98 154 100 164
rect 108 154 110 167
rect 128 147 130 161
rect 138 152 140 160
rect 148 150 150 158
rect 181 153 183 167
rect 192 147 194 167
rect 199 147 201 167
rect 219 147 221 161
rect 229 147 231 161
rect 239 154 241 164
rect 249 154 251 167
rect 281 154 283 167
rect 291 154 293 164
rect 301 147 303 161
rect 311 147 313 161
rect 331 147 333 167
rect 338 147 340 167
rect 349 153 351 167
rect 382 147 384 161
rect 392 152 394 160
rect 402 150 404 158
rect 435 153 437 167
rect 446 147 448 167
rect 453 147 455 167
rect 473 147 475 161
rect 483 147 485 161
rect 493 154 495 164
rect 503 154 505 167
rect 536 153 538 167
rect 547 147 549 167
rect 554 147 556 167
rect 574 147 576 161
rect 584 147 586 161
rect 594 154 596 164
rect 604 154 606 167
rect 635 153 637 167
rect 646 147 648 167
rect 653 147 655 167
rect 673 147 675 161
rect 683 147 685 161
rect 693 154 695 164
rect 703 154 705 167
rect 38 41 40 55
rect 48 42 50 50
rect 58 44 60 52
rect 79 35 81 49
rect 90 35 92 55
rect 97 35 99 55
rect 117 41 119 55
rect 127 41 129 55
rect 137 38 139 48
rect 147 35 149 48
rect 180 35 182 49
rect 191 35 193 55
rect 198 35 200 55
rect 218 41 220 55
rect 228 41 230 55
rect 238 38 240 48
rect 248 35 250 48
rect 281 35 283 49
rect 292 35 294 55
rect 299 35 301 55
rect 319 41 321 55
rect 329 41 331 55
rect 339 38 341 48
rect 349 35 351 48
rect 381 41 383 55
rect 391 42 393 50
rect 401 44 403 52
rect 434 35 436 49
rect 445 35 447 55
rect 452 35 454 55
rect 472 41 474 55
rect 482 41 484 55
rect 492 38 494 48
rect 502 35 504 48
rect 535 35 537 49
rect 546 35 548 55
rect 553 35 555 55
rect 573 41 575 55
rect 583 41 585 55
rect 593 38 595 48
rect 603 35 605 48
rect 634 35 636 49
rect 645 35 647 55
rect 652 35 654 55
rect 672 41 674 55
rect 682 41 684 55
rect 692 38 694 48
rect 702 35 704 48
<< pmos >>
rect 38 364 40 383
rect 48 364 50 383
rect 58 355 60 383
rect 78 364 80 383
rect 88 364 90 383
rect 98 355 100 383
rect 119 355 121 383
rect 129 355 131 383
rect 139 355 141 383
rect 157 355 159 380
rect 164 355 166 380
rect 174 358 176 371
rect 187 358 189 383
rect 215 358 217 383
rect 228 358 230 371
rect 238 355 240 380
rect 245 355 247 380
rect 263 355 265 383
rect 273 355 275 383
rect 283 355 285 383
rect 304 355 306 383
rect 314 364 316 383
rect 324 364 326 383
rect 344 355 346 383
rect 354 364 356 383
rect 364 364 366 383
rect 385 358 387 383
rect 398 358 400 371
rect 408 355 410 380
rect 415 355 417 380
rect 433 355 435 383
rect 443 355 445 383
rect 453 355 455 383
rect 474 355 476 383
rect 484 364 486 383
rect 494 364 496 383
rect 514 355 516 383
rect 524 364 526 383
rect 534 364 536 383
rect 554 364 556 383
rect 564 364 566 383
rect 574 355 576 383
rect 594 364 596 383
rect 604 364 606 383
rect 614 355 616 383
rect 635 355 637 383
rect 645 355 647 383
rect 655 355 657 383
rect 673 355 675 380
rect 680 355 682 380
rect 690 358 692 371
rect 703 358 705 383
rect 38 251 40 270
rect 48 251 50 270
rect 58 251 60 279
rect 78 251 80 270
rect 88 251 90 270
rect 98 251 100 279
rect 119 251 121 279
rect 129 251 131 279
rect 139 251 141 279
rect 157 254 159 279
rect 164 254 166 279
rect 174 263 176 276
rect 187 251 189 276
rect 215 251 217 276
rect 228 263 230 276
rect 238 254 240 279
rect 245 254 247 279
rect 263 251 265 279
rect 273 251 275 279
rect 283 251 285 279
rect 304 251 306 279
rect 314 251 316 270
rect 324 251 326 270
rect 344 251 346 279
rect 354 251 356 270
rect 364 251 366 270
rect 385 251 387 276
rect 398 263 400 276
rect 408 254 410 279
rect 415 254 417 279
rect 433 251 435 279
rect 443 251 445 279
rect 453 251 455 279
rect 474 251 476 279
rect 484 251 486 270
rect 494 251 496 270
rect 514 251 516 279
rect 524 251 526 270
rect 534 251 536 270
rect 554 251 556 270
rect 564 251 566 270
rect 574 251 576 279
rect 594 251 596 270
rect 604 251 606 270
rect 614 251 616 279
rect 635 251 637 279
rect 645 251 647 279
rect 655 251 657 279
rect 673 254 675 279
rect 680 254 682 279
rect 690 263 692 276
rect 703 251 705 276
rect 38 211 40 239
rect 51 211 53 239
rect 58 211 60 239
rect 79 211 81 239
rect 89 211 91 239
rect 99 211 101 239
rect 117 211 119 236
rect 124 211 126 236
rect 134 214 136 227
rect 147 214 149 239
rect 180 211 182 239
rect 190 211 192 239
rect 200 211 202 239
rect 218 211 220 236
rect 225 211 227 236
rect 235 214 237 227
rect 248 214 250 239
rect 282 211 284 239
rect 292 211 294 239
rect 302 211 304 239
rect 320 211 322 236
rect 327 211 329 236
rect 337 214 339 227
rect 350 214 352 239
rect 382 211 384 239
rect 395 211 397 239
rect 402 211 404 239
rect 435 211 437 239
rect 445 211 447 239
rect 455 211 457 239
rect 473 211 475 236
rect 480 211 482 236
rect 490 214 492 227
rect 503 214 505 239
rect 536 211 538 239
rect 546 211 548 239
rect 556 211 558 239
rect 574 211 576 236
rect 581 211 583 236
rect 591 214 593 227
rect 604 214 606 239
rect 635 211 637 239
rect 645 211 647 239
rect 655 211 657 239
rect 673 211 675 236
rect 680 211 682 236
rect 690 214 692 227
rect 703 214 705 239
rect 40 107 42 135
rect 50 107 52 135
rect 60 107 62 135
rect 78 110 80 135
rect 85 110 87 135
rect 95 119 97 132
rect 108 107 110 132
rect 128 107 130 135
rect 141 107 143 135
rect 148 107 150 135
rect 181 107 183 135
rect 191 107 193 135
rect 201 107 203 135
rect 219 110 221 135
rect 226 110 228 135
rect 236 119 238 132
rect 249 107 251 132
rect 281 107 283 132
rect 294 119 296 132
rect 304 110 306 135
rect 311 110 313 135
rect 329 107 331 135
rect 339 107 341 135
rect 349 107 351 135
rect 382 107 384 135
rect 395 107 397 135
rect 402 107 404 135
rect 435 107 437 135
rect 445 107 447 135
rect 455 107 457 135
rect 473 110 475 135
rect 480 110 482 135
rect 490 119 492 132
rect 503 107 505 132
rect 536 107 538 135
rect 546 107 548 135
rect 556 107 558 135
rect 574 110 576 135
rect 581 110 583 135
rect 591 119 593 132
rect 604 107 606 132
rect 635 107 637 135
rect 645 107 647 135
rect 655 107 657 135
rect 673 110 675 135
rect 680 110 682 135
rect 690 119 692 132
rect 703 107 705 132
rect 38 67 40 95
rect 51 67 53 95
rect 58 67 60 95
rect 79 67 81 95
rect 89 67 91 95
rect 99 67 101 95
rect 117 67 119 92
rect 124 67 126 92
rect 134 70 136 83
rect 147 70 149 95
rect 180 67 182 95
rect 190 67 192 95
rect 200 67 202 95
rect 218 67 220 92
rect 225 67 227 92
rect 235 70 237 83
rect 248 70 250 95
rect 281 67 283 95
rect 291 67 293 95
rect 301 67 303 95
rect 319 67 321 92
rect 326 67 328 92
rect 336 70 338 83
rect 349 70 351 95
rect 381 67 383 95
rect 394 67 396 95
rect 401 67 403 95
rect 434 67 436 95
rect 444 67 446 95
rect 454 67 456 95
rect 472 67 474 92
rect 479 67 481 92
rect 489 70 491 83
rect 502 70 504 95
rect 535 67 537 95
rect 545 67 547 95
rect 555 67 557 95
rect 573 67 575 92
rect 580 67 582 92
rect 590 70 592 83
rect 603 70 605 95
rect 634 67 636 95
rect 644 67 646 95
rect 654 67 656 95
rect 672 67 674 92
rect 679 67 681 92
rect 689 70 691 83
rect 702 70 704 95
<< polyct0 >>
rect 56 348 58 350
rect 96 348 98 350
rect 119 348 121 350
rect 129 348 131 350
rect 179 351 181 353
rect 185 341 187 343
rect 223 351 225 353
rect 217 341 219 343
rect 273 348 275 350
rect 283 348 285 350
rect 306 348 308 350
rect 346 348 348 350
rect 393 351 395 353
rect 387 341 389 343
rect 443 348 445 350
rect 453 348 455 350
rect 476 348 478 350
rect 516 348 518 350
rect 572 348 574 350
rect 612 348 614 350
rect 635 348 637 350
rect 645 348 647 350
rect 695 351 697 353
rect 701 341 703 343
rect 56 284 58 286
rect 96 284 98 286
rect 119 284 121 286
rect 129 284 131 286
rect 185 291 187 293
rect 179 281 181 283
rect 217 291 219 293
rect 223 281 225 283
rect 387 291 389 293
rect 273 284 275 286
rect 283 284 285 286
rect 306 284 308 286
rect 346 284 348 286
rect 393 281 395 283
rect 443 284 445 286
rect 453 284 455 286
rect 476 284 478 286
rect 516 284 518 286
rect 572 284 574 286
rect 612 284 614 286
rect 635 284 637 286
rect 645 284 647 286
rect 701 291 703 293
rect 695 281 697 283
rect 40 204 42 206
rect 79 204 81 206
rect 89 204 91 206
rect 139 207 141 209
rect 180 204 182 206
rect 190 204 192 206
rect 145 197 147 199
rect 240 207 242 209
rect 282 204 284 206
rect 292 204 294 206
rect 246 197 248 199
rect 342 207 344 209
rect 384 204 386 206
rect 435 204 437 206
rect 445 204 447 206
rect 348 197 350 199
rect 495 207 497 209
rect 536 204 538 206
rect 546 204 548 206
rect 501 197 503 199
rect 596 207 598 209
rect 635 204 637 206
rect 645 204 647 206
rect 602 197 604 199
rect 695 207 697 209
rect 701 197 703 199
rect 40 140 42 142
rect 50 140 52 142
rect 106 147 108 149
rect 100 137 102 139
rect 130 140 132 142
rect 181 140 183 142
rect 191 140 193 142
rect 247 147 249 149
rect 241 137 243 139
rect 283 147 285 149
rect 289 137 291 139
rect 339 140 341 142
rect 349 140 351 142
rect 384 140 386 142
rect 435 140 437 142
rect 445 140 447 142
rect 501 147 503 149
rect 495 137 497 139
rect 536 140 538 142
rect 546 140 548 142
rect 602 147 604 149
rect 596 137 598 139
rect 635 140 637 142
rect 645 140 647 142
rect 701 147 703 149
rect 695 137 697 139
rect 40 60 42 62
rect 79 60 81 62
rect 89 60 91 62
rect 139 63 141 65
rect 180 60 182 62
rect 190 60 192 62
rect 145 53 147 55
rect 240 63 242 65
rect 281 60 283 62
rect 291 60 293 62
rect 246 53 248 55
rect 341 63 343 65
rect 383 60 385 62
rect 434 60 436 62
rect 444 60 446 62
rect 347 53 349 55
rect 494 63 496 65
rect 535 60 537 62
rect 545 60 547 62
rect 500 53 502 55
rect 595 63 597 65
rect 634 60 636 62
rect 644 60 646 62
rect 601 53 603 55
rect 694 63 696 65
rect 700 53 702 55
<< polyct1 >>
rect 36 356 38 358
rect 76 356 78 358
rect 46 348 48 350
rect 86 348 88 350
rect 139 348 141 350
rect 146 348 148 350
rect 165 348 167 350
rect 326 356 328 358
rect 237 348 239 350
rect 256 348 258 350
rect 263 348 265 350
rect 316 348 318 350
rect 366 356 368 358
rect 356 348 358 350
rect 496 356 498 358
rect 407 348 409 350
rect 426 348 428 350
rect 433 348 435 350
rect 486 348 488 350
rect 536 356 538 358
rect 552 356 554 358
rect 526 348 528 350
rect 592 356 594 358
rect 562 348 564 350
rect 602 348 604 350
rect 655 348 657 350
rect 662 348 664 350
rect 681 348 683 350
rect 46 284 48 286
rect 36 276 38 278
rect 86 284 88 286
rect 139 284 141 286
rect 146 284 148 286
rect 165 284 167 286
rect 76 276 78 278
rect 237 284 239 286
rect 256 284 258 286
rect 263 284 265 286
rect 316 284 318 286
rect 356 284 358 286
rect 326 276 328 278
rect 366 276 368 278
rect 407 284 409 286
rect 426 284 428 286
rect 433 284 435 286
rect 486 284 488 286
rect 526 284 528 286
rect 496 276 498 278
rect 562 284 564 286
rect 536 276 538 278
rect 552 276 554 278
rect 602 284 604 286
rect 655 284 657 286
rect 662 284 664 286
rect 681 284 683 286
rect 592 276 594 278
rect 50 204 52 206
rect 63 204 65 206
rect 99 204 101 206
rect 106 204 108 206
rect 125 204 127 206
rect 200 204 202 206
rect 207 204 209 206
rect 226 204 228 206
rect 302 204 304 206
rect 309 204 311 206
rect 328 204 330 206
rect 394 204 396 206
rect 407 204 409 206
rect 455 204 457 206
rect 462 204 464 206
rect 481 204 483 206
rect 556 204 558 206
rect 563 204 565 206
rect 582 204 584 206
rect 655 204 657 206
rect 662 204 664 206
rect 681 204 683 206
rect 60 140 62 142
rect 67 140 69 142
rect 86 140 88 142
rect 140 140 142 142
rect 153 140 155 142
rect 201 140 203 142
rect 208 140 210 142
rect 227 140 229 142
rect 303 140 305 142
rect 322 140 324 142
rect 329 140 331 142
rect 394 140 396 142
rect 407 140 409 142
rect 455 140 457 142
rect 462 140 464 142
rect 481 140 483 142
rect 556 140 558 142
rect 563 140 565 142
rect 582 140 584 142
rect 655 140 657 142
rect 662 140 664 142
rect 681 140 683 142
rect 50 60 52 62
rect 63 60 65 62
rect 99 60 101 62
rect 106 60 108 62
rect 125 60 127 62
rect 200 60 202 62
rect 207 60 209 62
rect 226 60 228 62
rect 301 60 303 62
rect 308 60 310 62
rect 327 60 329 62
rect 393 60 395 62
rect 406 60 408 62
rect 454 60 456 62
rect 461 60 463 62
rect 480 60 482 62
rect 555 60 557 62
rect 562 60 564 62
rect 581 60 583 62
rect 654 60 656 62
rect 661 60 663 62
rect 680 60 682 62
<< ndifct0 >>
rect 33 332 35 334
rect 73 332 75 334
rect 125 325 127 327
rect 152 339 154 341
rect 142 332 144 334
rect 152 332 154 334
rect 162 339 164 341
rect 172 331 174 333
rect 182 328 184 330
rect 220 328 222 330
rect 230 331 232 333
rect 240 339 242 341
rect 250 339 252 341
rect 250 332 252 334
rect 260 332 262 334
rect 277 325 279 327
rect 329 332 331 334
rect 369 332 371 334
rect 390 328 392 330
rect 400 331 402 333
rect 410 339 412 341
rect 420 339 422 341
rect 420 332 422 334
rect 430 332 432 334
rect 447 325 449 327
rect 499 332 501 334
rect 539 332 541 334
rect 549 332 551 334
rect 589 332 591 334
rect 641 325 643 327
rect 668 339 670 341
rect 658 332 660 334
rect 668 332 670 334
rect 678 339 680 341
rect 688 331 690 333
rect 698 328 700 330
rect 33 300 35 302
rect 73 300 75 302
rect 125 307 127 309
rect 142 300 144 302
rect 152 300 154 302
rect 152 293 154 295
rect 162 293 164 295
rect 172 301 174 303
rect 182 304 184 306
rect 220 304 222 306
rect 230 301 232 303
rect 240 293 242 295
rect 250 300 252 302
rect 260 300 262 302
rect 250 293 252 295
rect 277 307 279 309
rect 329 300 331 302
rect 369 300 371 302
rect 390 304 392 306
rect 400 301 402 303
rect 410 293 412 295
rect 420 300 422 302
rect 430 300 432 302
rect 420 293 422 295
rect 447 307 449 309
rect 499 300 501 302
rect 539 300 541 302
rect 549 300 551 302
rect 589 300 591 302
rect 641 307 643 309
rect 658 300 660 302
rect 668 300 670 302
rect 668 293 670 295
rect 678 293 680 295
rect 688 301 690 303
rect 698 304 700 306
rect 43 188 45 190
rect 53 190 55 192
rect 63 190 65 192
rect 85 181 87 183
rect 112 195 114 197
rect 102 188 104 190
rect 112 188 114 190
rect 122 195 124 197
rect 132 187 134 189
rect 142 184 144 186
rect 186 181 188 183
rect 213 195 215 197
rect 203 188 205 190
rect 213 188 215 190
rect 223 195 225 197
rect 233 187 235 189
rect 243 184 245 186
rect 288 181 290 183
rect 315 195 317 197
rect 305 188 307 190
rect 315 188 317 190
rect 325 195 327 197
rect 335 187 337 189
rect 345 184 347 186
rect 387 188 389 190
rect 397 190 399 192
rect 407 190 409 192
rect 441 181 443 183
rect 468 195 470 197
rect 458 188 460 190
rect 468 188 470 190
rect 478 195 480 197
rect 488 187 490 189
rect 498 184 500 186
rect 542 181 544 183
rect 569 195 571 197
rect 559 188 561 190
rect 569 188 571 190
rect 579 195 581 197
rect 589 187 591 189
rect 599 184 601 186
rect 641 181 643 183
rect 668 195 670 197
rect 658 188 660 190
rect 668 188 670 190
rect 678 195 680 197
rect 688 187 690 189
rect 698 184 700 186
rect 46 163 48 165
rect 63 156 65 158
rect 73 156 75 158
rect 73 149 75 151
rect 83 149 85 151
rect 93 157 95 159
rect 103 160 105 162
rect 133 156 135 158
rect 143 154 145 156
rect 153 154 155 156
rect 187 163 189 165
rect 204 156 206 158
rect 214 156 216 158
rect 214 149 216 151
rect 224 149 226 151
rect 234 157 236 159
rect 244 160 246 162
rect 286 160 288 162
rect 296 157 298 159
rect 306 149 308 151
rect 316 156 318 158
rect 326 156 328 158
rect 316 149 318 151
rect 343 163 345 165
rect 387 156 389 158
rect 397 154 399 156
rect 407 154 409 156
rect 441 163 443 165
rect 458 156 460 158
rect 468 156 470 158
rect 468 149 470 151
rect 478 149 480 151
rect 488 157 490 159
rect 498 160 500 162
rect 542 163 544 165
rect 559 156 561 158
rect 569 156 571 158
rect 569 149 571 151
rect 579 149 581 151
rect 589 157 591 159
rect 599 160 601 162
rect 641 163 643 165
rect 658 156 660 158
rect 668 156 670 158
rect 668 149 670 151
rect 678 149 680 151
rect 688 157 690 159
rect 698 160 700 162
rect 43 44 45 46
rect 53 46 55 48
rect 63 46 65 48
rect 85 37 87 39
rect 112 51 114 53
rect 102 44 104 46
rect 112 44 114 46
rect 122 51 124 53
rect 132 43 134 45
rect 142 40 144 42
rect 186 37 188 39
rect 213 51 215 53
rect 203 44 205 46
rect 213 44 215 46
rect 223 51 225 53
rect 233 43 235 45
rect 243 40 245 42
rect 287 37 289 39
rect 314 51 316 53
rect 304 44 306 46
rect 314 44 316 46
rect 324 51 326 53
rect 334 43 336 45
rect 344 40 346 42
rect 386 44 388 46
rect 396 46 398 48
rect 406 46 408 48
rect 440 37 442 39
rect 467 51 469 53
rect 457 44 459 46
rect 467 44 469 46
rect 477 51 479 53
rect 487 43 489 45
rect 497 40 499 42
rect 541 37 543 39
rect 568 51 570 53
rect 558 44 560 46
rect 568 44 570 46
rect 578 51 580 53
rect 588 43 590 45
rect 598 40 600 42
rect 640 37 642 39
rect 667 51 669 53
rect 657 44 659 46
rect 667 44 669 46
rect 677 51 679 53
rect 687 43 689 45
rect 697 40 699 42
<< ndifct1 >>
rect 63 339 65 341
rect 63 331 65 333
rect 103 339 105 341
rect 103 331 105 333
rect 114 332 116 334
rect 52 322 54 324
rect 92 322 94 324
rect 192 332 194 334
rect 210 332 212 334
rect 299 339 301 341
rect 288 332 290 334
rect 299 331 301 333
rect 339 339 341 341
rect 339 331 341 333
rect 380 332 382 334
rect 310 322 312 324
rect 350 322 352 324
rect 469 339 471 341
rect 458 332 460 334
rect 469 331 471 333
rect 509 339 511 341
rect 509 331 511 333
rect 579 339 581 341
rect 579 331 581 333
rect 480 322 482 324
rect 520 322 522 324
rect 619 339 621 341
rect 619 331 621 333
rect 630 332 632 334
rect 568 322 570 324
rect 608 322 610 324
rect 708 332 710 334
rect 52 310 54 312
rect 92 310 94 312
rect 63 301 65 303
rect 63 293 65 295
rect 103 301 105 303
rect 114 300 116 302
rect 103 293 105 295
rect 192 300 194 302
rect 210 300 212 302
rect 310 310 312 312
rect 350 310 352 312
rect 288 300 290 302
rect 299 301 301 303
rect 299 293 301 295
rect 339 301 341 303
rect 339 293 341 295
rect 380 300 382 302
rect 480 310 482 312
rect 520 310 522 312
rect 458 300 460 302
rect 469 301 471 303
rect 469 293 471 295
rect 568 310 570 312
rect 608 310 610 312
rect 509 301 511 303
rect 509 293 511 295
rect 579 301 581 303
rect 579 293 581 295
rect 619 301 621 303
rect 630 300 632 302
rect 619 293 621 295
rect 708 300 710 302
rect 33 195 35 197
rect 33 188 35 190
rect 74 188 76 190
rect 152 188 154 190
rect 175 188 177 190
rect 253 188 255 190
rect 277 188 279 190
rect 377 195 379 197
rect 355 188 357 190
rect 377 188 379 190
rect 430 188 432 190
rect 508 188 510 190
rect 531 188 533 190
rect 609 188 611 190
rect 630 188 632 190
rect 708 188 710 190
rect 35 156 37 158
rect 113 156 115 158
rect 123 156 125 158
rect 123 149 125 151
rect 176 156 178 158
rect 254 156 256 158
rect 276 156 278 158
rect 354 156 356 158
rect 377 156 379 158
rect 377 149 379 151
rect 430 156 432 158
rect 508 156 510 158
rect 531 156 533 158
rect 609 156 611 158
rect 630 156 632 158
rect 708 156 710 158
rect 33 51 35 53
rect 33 44 35 46
rect 74 44 76 46
rect 152 44 154 46
rect 175 44 177 46
rect 253 44 255 46
rect 276 44 278 46
rect 376 51 378 53
rect 354 44 356 46
rect 376 44 378 46
rect 429 44 431 46
rect 507 44 509 46
rect 530 44 532 46
rect 608 44 610 46
rect 629 44 631 46
rect 707 44 709 46
<< ptiect1 >>
rect 404 178 406 180
rect 150 166 152 168
rect 404 166 406 168
rect 60 34 62 36
rect 403 34 405 36
<< pdifct0 >>
rect 33 379 35 381
rect 33 372 35 374
rect 43 373 45 375
rect 43 366 45 368
rect 53 379 55 381
rect 53 372 55 374
rect 73 379 75 381
rect 73 372 75 374
rect 83 373 85 375
rect 83 366 85 368
rect 93 379 95 381
rect 93 372 95 374
rect 124 379 126 381
rect 124 372 126 374
rect 134 371 136 373
rect 134 364 136 366
rect 146 379 148 381
rect 146 372 148 374
rect 181 379 183 381
rect 169 360 171 362
rect 221 379 223 381
rect 233 360 235 362
rect 256 379 258 381
rect 256 372 258 374
rect 268 371 270 373
rect 268 364 270 366
rect 278 379 280 381
rect 278 372 280 374
rect 309 379 311 381
rect 309 372 311 374
rect 319 373 321 375
rect 319 366 321 368
rect 329 379 331 381
rect 329 372 331 374
rect 349 379 351 381
rect 349 372 351 374
rect 359 373 361 375
rect 359 366 361 368
rect 369 379 371 381
rect 369 372 371 374
rect 391 379 393 381
rect 403 360 405 362
rect 426 379 428 381
rect 426 372 428 374
rect 438 371 440 373
rect 438 364 440 366
rect 448 379 450 381
rect 448 372 450 374
rect 479 379 481 381
rect 479 372 481 374
rect 489 373 491 375
rect 489 366 491 368
rect 499 379 501 381
rect 499 372 501 374
rect 519 379 521 381
rect 519 372 521 374
rect 529 373 531 375
rect 529 366 531 368
rect 539 379 541 381
rect 539 372 541 374
rect 549 379 551 381
rect 549 372 551 374
rect 559 373 561 375
rect 559 366 561 368
rect 569 379 571 381
rect 569 372 571 374
rect 589 379 591 381
rect 589 372 591 374
rect 599 373 601 375
rect 599 366 601 368
rect 609 379 611 381
rect 609 372 611 374
rect 640 379 642 381
rect 640 372 642 374
rect 650 371 652 373
rect 650 364 652 366
rect 662 379 664 381
rect 662 372 664 374
rect 697 379 699 381
rect 685 360 687 362
rect 33 260 35 262
rect 33 253 35 255
rect 43 266 45 268
rect 43 259 45 261
rect 53 260 55 262
rect 53 253 55 255
rect 73 260 75 262
rect 73 253 75 255
rect 83 266 85 268
rect 83 259 85 261
rect 93 260 95 262
rect 93 253 95 255
rect 124 260 126 262
rect 124 253 126 255
rect 134 268 136 270
rect 134 261 136 263
rect 146 260 148 262
rect 146 253 148 255
rect 169 272 171 274
rect 181 253 183 255
rect 233 272 235 274
rect 221 253 223 255
rect 256 260 258 262
rect 256 253 258 255
rect 268 268 270 270
rect 268 261 270 263
rect 278 260 280 262
rect 278 253 280 255
rect 309 260 311 262
rect 309 253 311 255
rect 319 266 321 268
rect 319 259 321 261
rect 329 260 331 262
rect 329 253 331 255
rect 349 260 351 262
rect 349 253 351 255
rect 359 266 361 268
rect 359 259 361 261
rect 369 260 371 262
rect 369 253 371 255
rect 403 272 405 274
rect 391 253 393 255
rect 426 260 428 262
rect 426 253 428 255
rect 438 268 440 270
rect 438 261 440 263
rect 448 260 450 262
rect 448 253 450 255
rect 479 260 481 262
rect 479 253 481 255
rect 489 266 491 268
rect 489 259 491 261
rect 499 260 501 262
rect 499 253 501 255
rect 519 260 521 262
rect 519 253 521 255
rect 529 266 531 268
rect 529 259 531 261
rect 539 260 541 262
rect 539 253 541 255
rect 549 260 551 262
rect 549 253 551 255
rect 559 266 561 268
rect 559 259 561 261
rect 569 260 571 262
rect 569 253 571 255
rect 589 260 591 262
rect 589 253 591 255
rect 599 266 601 268
rect 599 259 601 261
rect 609 260 611 262
rect 609 253 611 255
rect 640 260 642 262
rect 640 253 642 255
rect 650 268 652 270
rect 650 261 652 263
rect 662 260 664 262
rect 662 253 664 255
rect 685 272 687 274
rect 697 253 699 255
rect 63 229 65 231
rect 84 235 86 237
rect 84 228 86 230
rect 94 227 96 229
rect 94 220 96 222
rect 106 235 108 237
rect 106 228 108 230
rect 141 235 143 237
rect 129 216 131 218
rect 185 235 187 237
rect 185 228 187 230
rect 195 227 197 229
rect 195 220 197 222
rect 207 235 209 237
rect 207 228 209 230
rect 242 235 244 237
rect 230 216 232 218
rect 287 235 289 237
rect 287 228 289 230
rect 297 227 299 229
rect 297 220 299 222
rect 309 235 311 237
rect 309 228 311 230
rect 344 235 346 237
rect 332 216 334 218
rect 407 229 409 231
rect 440 235 442 237
rect 440 228 442 230
rect 450 227 452 229
rect 450 220 452 222
rect 462 235 464 237
rect 462 228 464 230
rect 497 235 499 237
rect 485 216 487 218
rect 541 235 543 237
rect 541 228 543 230
rect 551 227 553 229
rect 551 220 553 222
rect 563 235 565 237
rect 563 228 565 230
rect 598 235 600 237
rect 586 216 588 218
rect 640 235 642 237
rect 640 228 642 230
rect 650 227 652 229
rect 650 220 652 222
rect 662 235 664 237
rect 662 228 664 230
rect 697 235 699 237
rect 685 216 687 218
rect 45 116 47 118
rect 45 109 47 111
rect 55 124 57 126
rect 55 117 57 119
rect 67 116 69 118
rect 67 109 69 111
rect 90 128 92 130
rect 102 109 104 111
rect 153 115 155 117
rect 186 116 188 118
rect 186 109 188 111
rect 196 124 198 126
rect 196 117 198 119
rect 208 116 210 118
rect 208 109 210 111
rect 231 128 233 130
rect 243 109 245 111
rect 299 128 301 130
rect 287 109 289 111
rect 322 116 324 118
rect 322 109 324 111
rect 334 124 336 126
rect 334 117 336 119
rect 344 116 346 118
rect 344 109 346 111
rect 407 115 409 117
rect 440 116 442 118
rect 440 109 442 111
rect 450 124 452 126
rect 450 117 452 119
rect 462 116 464 118
rect 462 109 464 111
rect 485 128 487 130
rect 497 109 499 111
rect 541 116 543 118
rect 541 109 543 111
rect 551 124 553 126
rect 551 117 553 119
rect 563 116 565 118
rect 563 109 565 111
rect 586 128 588 130
rect 598 109 600 111
rect 640 116 642 118
rect 640 109 642 111
rect 650 124 652 126
rect 650 117 652 119
rect 662 116 664 118
rect 662 109 664 111
rect 685 128 687 130
rect 697 109 699 111
rect 63 85 65 87
rect 84 91 86 93
rect 84 84 86 86
rect 94 83 96 85
rect 94 76 96 78
rect 106 91 108 93
rect 106 84 108 86
rect 141 91 143 93
rect 129 72 131 74
rect 185 91 187 93
rect 185 84 187 86
rect 195 83 197 85
rect 195 76 197 78
rect 207 91 209 93
rect 207 84 209 86
rect 242 91 244 93
rect 230 72 232 74
rect 286 91 288 93
rect 286 84 288 86
rect 296 83 298 85
rect 296 76 298 78
rect 308 91 310 93
rect 308 84 310 86
rect 343 91 345 93
rect 331 72 333 74
rect 406 85 408 87
rect 439 91 441 93
rect 439 84 441 86
rect 449 83 451 85
rect 449 76 451 78
rect 461 91 463 93
rect 461 84 463 86
rect 496 91 498 93
rect 484 72 486 74
rect 540 91 542 93
rect 540 84 542 86
rect 550 83 552 85
rect 550 76 552 78
rect 562 91 564 93
rect 562 84 564 86
rect 597 91 599 93
rect 585 72 587 74
rect 639 91 641 93
rect 639 84 641 86
rect 649 83 651 85
rect 649 76 651 78
rect 661 91 663 93
rect 661 84 663 86
rect 696 91 698 93
rect 684 72 686 74
<< pdifct1 >>
rect 63 372 65 374
rect 63 365 65 367
rect 103 372 105 374
rect 103 365 105 367
rect 114 364 116 366
rect 114 357 116 359
rect 192 367 194 369
rect 192 360 194 362
rect 210 367 212 369
rect 210 360 212 362
rect 299 372 301 374
rect 288 364 290 366
rect 299 365 301 367
rect 288 357 290 359
rect 339 372 341 374
rect 339 365 341 367
rect 380 367 382 369
rect 380 360 382 362
rect 469 372 471 374
rect 458 364 460 366
rect 469 365 471 367
rect 458 357 460 359
rect 509 372 511 374
rect 509 365 511 367
rect 579 372 581 374
rect 579 365 581 367
rect 619 372 621 374
rect 619 365 621 367
rect 630 364 632 366
rect 630 357 632 359
rect 708 367 710 369
rect 708 360 710 362
rect 63 267 65 269
rect 63 260 65 262
rect 114 275 116 277
rect 103 267 105 269
rect 103 260 105 262
rect 192 272 194 274
rect 192 265 194 267
rect 210 272 212 274
rect 210 265 212 267
rect 288 275 290 277
rect 288 268 290 270
rect 299 267 301 269
rect 299 260 301 262
rect 339 267 341 269
rect 339 260 341 262
rect 380 272 382 274
rect 380 265 382 267
rect 458 275 460 277
rect 458 268 460 270
rect 469 267 471 269
rect 469 260 471 262
rect 509 267 511 269
rect 509 260 511 262
rect 579 267 581 269
rect 579 260 581 262
rect 630 275 632 277
rect 619 267 621 269
rect 630 268 632 270
rect 619 260 621 262
rect 708 272 710 274
rect 708 265 710 267
rect 33 229 35 231
rect 33 222 35 224
rect 44 238 46 240
rect 74 220 76 222
rect 74 213 76 215
rect 152 223 154 225
rect 152 216 154 218
rect 175 220 177 222
rect 175 213 177 215
rect 253 223 255 225
rect 253 216 255 218
rect 277 220 279 222
rect 277 213 279 215
rect 377 229 379 231
rect 355 223 357 225
rect 377 222 379 224
rect 355 216 357 218
rect 388 238 390 240
rect 430 220 432 222
rect 430 213 432 215
rect 508 223 510 225
rect 508 216 510 218
rect 531 220 533 222
rect 531 213 533 215
rect 609 223 611 225
rect 609 216 611 218
rect 630 220 632 222
rect 630 213 632 215
rect 708 223 710 225
rect 708 216 710 218
rect 35 131 37 133
rect 35 124 37 126
rect 113 128 115 130
rect 113 121 115 123
rect 123 122 125 124
rect 123 115 125 117
rect 134 106 136 108
rect 176 131 178 133
rect 176 124 178 126
rect 254 128 256 130
rect 254 121 256 123
rect 276 128 278 130
rect 276 121 278 123
rect 354 131 356 133
rect 354 124 356 126
rect 377 122 379 124
rect 377 115 379 117
rect 388 106 390 108
rect 430 131 432 133
rect 430 124 432 126
rect 508 128 510 130
rect 508 121 510 123
rect 531 131 533 133
rect 531 124 533 126
rect 609 128 611 130
rect 609 121 611 123
rect 630 131 632 133
rect 630 124 632 126
rect 708 128 710 130
rect 708 121 710 123
rect 33 85 35 87
rect 33 78 35 80
rect 44 94 46 96
rect 74 76 76 78
rect 74 69 76 71
rect 152 79 154 81
rect 152 72 154 74
rect 175 76 177 78
rect 175 69 177 71
rect 253 79 255 81
rect 253 72 255 74
rect 276 76 278 78
rect 276 69 278 71
rect 376 85 378 87
rect 354 79 356 81
rect 376 78 378 80
rect 354 72 356 74
rect 387 94 389 96
rect 429 76 431 78
rect 429 69 431 71
rect 507 79 509 81
rect 507 72 509 74
rect 530 76 532 78
rect 530 69 532 71
rect 608 79 610 81
rect 608 72 610 74
rect 629 76 631 78
rect 629 69 631 71
rect 707 79 709 81
rect 707 72 709 74
<< alu0 >>
rect 31 379 33 381
rect 35 379 37 381
rect 31 374 37 379
rect 51 379 53 381
rect 55 379 57 381
rect 31 372 33 374
rect 35 372 37 374
rect 31 371 37 372
rect 41 375 47 376
rect 41 373 43 375
rect 45 373 47 375
rect 41 368 47 373
rect 51 374 57 379
rect 71 379 73 381
rect 75 379 77 381
rect 51 372 53 374
rect 55 372 57 374
rect 51 371 57 372
rect 41 366 43 368
rect 45 367 47 368
rect 71 374 77 379
rect 91 379 93 381
rect 95 379 97 381
rect 71 372 73 374
rect 75 372 77 374
rect 71 371 77 372
rect 81 375 87 376
rect 81 373 83 375
rect 85 373 87 375
rect 81 368 87 373
rect 91 374 97 379
rect 122 379 124 381
rect 126 379 128 381
rect 91 372 93 374
rect 95 372 97 374
rect 91 371 97 372
rect 45 366 55 367
rect 41 363 55 366
rect 51 359 55 363
rect 51 355 59 359
rect 55 350 59 355
rect 55 348 56 350
rect 58 348 59 350
rect 55 343 59 348
rect 47 339 59 343
rect 47 335 51 339
rect 62 336 63 343
rect 81 366 83 368
rect 85 367 87 368
rect 122 374 128 379
rect 144 379 146 381
rect 148 379 150 381
rect 122 372 124 374
rect 126 372 128 374
rect 122 371 128 372
rect 133 373 137 375
rect 133 371 134 373
rect 136 371 137 373
rect 144 374 150 379
rect 179 379 181 381
rect 183 379 185 381
rect 179 378 185 379
rect 219 379 221 381
rect 223 379 225 381
rect 219 378 225 379
rect 254 379 256 381
rect 258 379 260 381
rect 144 372 146 374
rect 148 372 150 374
rect 144 371 150 372
rect 85 366 95 367
rect 81 363 95 366
rect 91 359 95 363
rect 91 355 99 359
rect 95 350 99 355
rect 95 348 96 350
rect 98 348 99 350
rect 95 343 99 348
rect 87 339 99 343
rect 31 334 51 335
rect 31 332 33 334
rect 35 332 51 334
rect 31 331 51 332
rect 87 335 91 339
rect 102 336 103 343
rect 71 334 91 335
rect 71 332 73 334
rect 75 332 91 334
rect 71 331 91 332
rect 133 367 137 371
rect 156 367 180 371
rect 120 366 160 367
rect 120 364 134 366
rect 136 364 160 366
rect 120 363 160 364
rect 120 352 124 363
rect 168 362 172 364
rect 176 363 182 367
rect 168 360 169 362
rect 171 360 172 362
rect 168 359 172 360
rect 168 355 175 359
rect 118 350 124 352
rect 118 348 119 350
rect 121 348 124 350
rect 118 346 124 348
rect 128 350 132 355
rect 128 348 129 350
rect 131 348 132 350
rect 128 346 132 348
rect 120 343 124 346
rect 120 339 140 343
rect 136 335 140 339
rect 171 344 175 355
rect 178 353 182 363
rect 178 351 179 353
rect 181 351 182 353
rect 178 349 182 351
rect 171 343 189 344
rect 151 341 155 343
rect 171 342 185 343
rect 151 339 152 341
rect 154 339 155 341
rect 136 334 146 335
rect 136 332 142 334
rect 144 332 146 334
rect 136 331 146 332
rect 151 334 155 339
rect 160 341 185 342
rect 187 341 189 343
rect 160 339 162 341
rect 164 340 189 341
rect 164 339 175 340
rect 160 338 175 339
rect 151 332 152 334
rect 154 333 176 334
rect 154 332 172 333
rect 151 331 172 332
rect 174 331 176 333
rect 151 330 176 331
rect 181 330 185 332
rect 254 374 260 379
rect 276 379 278 381
rect 280 379 282 381
rect 254 372 256 374
rect 258 372 260 374
rect 254 371 260 372
rect 267 373 271 375
rect 267 371 268 373
rect 270 371 271 373
rect 276 374 282 379
rect 307 379 309 381
rect 311 379 313 381
rect 276 372 278 374
rect 280 372 282 374
rect 276 371 282 372
rect 224 367 248 371
rect 267 367 271 371
rect 222 363 228 367
rect 244 366 284 367
rect 244 364 268 366
rect 270 364 284 366
rect 222 353 226 363
rect 232 362 236 364
rect 244 363 284 364
rect 232 360 233 362
rect 235 360 236 362
rect 232 359 236 360
rect 222 351 223 353
rect 225 351 226 353
rect 222 349 226 351
rect 229 355 236 359
rect 229 344 233 355
rect 272 350 276 355
rect 272 348 273 350
rect 275 348 276 350
rect 215 343 233 344
rect 215 341 217 343
rect 219 342 233 343
rect 219 341 244 342
rect 215 340 240 341
rect 229 339 240 340
rect 242 339 244 341
rect 229 338 244 339
rect 249 341 253 343
rect 249 339 250 341
rect 252 339 253 341
rect 249 334 253 339
rect 272 346 276 348
rect 280 352 284 363
rect 280 350 286 352
rect 280 348 283 350
rect 285 348 286 350
rect 280 346 286 348
rect 280 343 284 346
rect 264 339 284 343
rect 264 335 268 339
rect 228 333 250 334
rect 219 330 223 332
rect 228 331 230 333
rect 232 332 250 333
rect 252 332 253 334
rect 232 331 253 332
rect 258 334 268 335
rect 258 332 260 334
rect 262 332 268 334
rect 258 331 268 332
rect 307 374 313 379
rect 327 379 329 381
rect 331 379 333 381
rect 307 372 309 374
rect 311 372 313 374
rect 307 371 313 372
rect 317 375 323 376
rect 317 373 319 375
rect 321 373 323 375
rect 317 368 323 373
rect 327 374 333 379
rect 347 379 349 381
rect 351 379 353 381
rect 327 372 329 374
rect 331 372 333 374
rect 327 371 333 372
rect 317 367 319 368
rect 309 366 319 367
rect 321 366 323 368
rect 309 363 323 366
rect 309 359 313 363
rect 305 355 313 359
rect 347 374 353 379
rect 367 379 369 381
rect 371 379 373 381
rect 347 372 349 374
rect 351 372 353 374
rect 347 371 353 372
rect 357 375 363 376
rect 357 373 359 375
rect 361 373 363 375
rect 357 368 363 373
rect 367 374 373 379
rect 389 379 391 381
rect 393 379 395 381
rect 389 378 395 379
rect 424 379 426 381
rect 428 379 430 381
rect 367 372 369 374
rect 371 372 373 374
rect 367 371 373 372
rect 424 374 430 379
rect 446 379 448 381
rect 450 379 452 381
rect 424 372 426 374
rect 428 372 430 374
rect 424 371 430 372
rect 437 373 441 375
rect 437 371 438 373
rect 440 371 441 373
rect 446 374 452 379
rect 477 379 479 381
rect 481 379 483 381
rect 446 372 448 374
rect 450 372 452 374
rect 446 371 452 372
rect 357 367 359 368
rect 349 366 359 367
rect 361 366 363 368
rect 349 363 363 366
rect 305 350 309 355
rect 305 348 306 350
rect 308 348 309 350
rect 305 343 309 348
rect 301 336 302 343
rect 305 339 317 343
rect 313 335 317 339
rect 349 359 353 363
rect 345 355 353 359
rect 394 367 418 371
rect 437 367 441 371
rect 392 363 398 367
rect 414 366 454 367
rect 414 364 438 366
rect 440 364 454 366
rect 345 350 349 355
rect 345 348 346 350
rect 348 348 349 350
rect 345 343 349 348
rect 341 336 342 343
rect 345 339 357 343
rect 313 334 333 335
rect 313 332 329 334
rect 331 332 333 334
rect 313 331 333 332
rect 353 335 357 339
rect 392 353 396 363
rect 402 362 406 364
rect 414 363 454 364
rect 402 360 403 362
rect 405 360 406 362
rect 402 359 406 360
rect 392 351 393 353
rect 395 351 396 353
rect 392 349 396 351
rect 399 355 406 359
rect 399 344 403 355
rect 442 350 446 355
rect 442 348 443 350
rect 445 348 446 350
rect 385 343 403 344
rect 385 341 387 343
rect 389 342 403 343
rect 389 341 414 342
rect 385 340 410 341
rect 399 339 410 340
rect 412 339 414 341
rect 399 338 414 339
rect 419 341 423 343
rect 419 339 420 341
rect 422 339 423 341
rect 353 334 373 335
rect 353 332 369 334
rect 371 332 373 334
rect 353 331 373 332
rect 419 334 423 339
rect 442 346 446 348
rect 450 352 454 363
rect 450 350 456 352
rect 450 348 453 350
rect 455 348 456 350
rect 450 346 456 348
rect 450 343 454 346
rect 434 339 454 343
rect 434 335 438 339
rect 398 333 420 334
rect 228 330 253 331
rect 389 330 393 332
rect 398 331 400 333
rect 402 332 420 333
rect 422 332 423 334
rect 402 331 423 332
rect 428 334 438 335
rect 428 332 430 334
rect 432 332 438 334
rect 428 331 438 332
rect 477 374 483 379
rect 497 379 499 381
rect 501 379 503 381
rect 477 372 479 374
rect 481 372 483 374
rect 477 371 483 372
rect 487 375 493 376
rect 487 373 489 375
rect 491 373 493 375
rect 487 368 493 373
rect 497 374 503 379
rect 517 379 519 381
rect 521 379 523 381
rect 497 372 499 374
rect 501 372 503 374
rect 497 371 503 372
rect 487 367 489 368
rect 479 366 489 367
rect 491 366 493 368
rect 479 363 493 366
rect 479 359 483 363
rect 475 355 483 359
rect 517 374 523 379
rect 537 379 539 381
rect 541 379 543 381
rect 517 372 519 374
rect 521 372 523 374
rect 517 371 523 372
rect 527 375 533 376
rect 527 373 529 375
rect 531 373 533 375
rect 527 368 533 373
rect 537 374 543 379
rect 537 372 539 374
rect 541 372 543 374
rect 537 371 543 372
rect 547 379 549 381
rect 551 379 553 381
rect 547 374 553 379
rect 567 379 569 381
rect 571 379 573 381
rect 547 372 549 374
rect 551 372 553 374
rect 547 371 553 372
rect 557 375 563 376
rect 557 373 559 375
rect 561 373 563 375
rect 557 368 563 373
rect 567 374 573 379
rect 587 379 589 381
rect 591 379 593 381
rect 567 372 569 374
rect 571 372 573 374
rect 567 371 573 372
rect 527 367 529 368
rect 519 366 529 367
rect 531 366 533 368
rect 519 363 533 366
rect 475 350 479 355
rect 475 348 476 350
rect 478 348 479 350
rect 475 343 479 348
rect 471 336 472 343
rect 475 339 487 343
rect 483 335 487 339
rect 519 359 523 363
rect 515 355 523 359
rect 557 366 559 368
rect 561 367 563 368
rect 587 374 593 379
rect 607 379 609 381
rect 611 379 613 381
rect 587 372 589 374
rect 591 372 593 374
rect 587 371 593 372
rect 597 375 603 376
rect 597 373 599 375
rect 601 373 603 375
rect 597 368 603 373
rect 607 374 613 379
rect 638 379 640 381
rect 642 379 644 381
rect 607 372 609 374
rect 611 372 613 374
rect 607 371 613 372
rect 561 366 571 367
rect 557 363 571 366
rect 567 359 571 363
rect 567 355 575 359
rect 515 350 519 355
rect 515 348 516 350
rect 518 348 519 350
rect 515 343 519 348
rect 511 336 512 343
rect 515 339 527 343
rect 483 334 503 335
rect 483 332 499 334
rect 501 332 503 334
rect 483 331 503 332
rect 523 335 527 339
rect 571 350 575 355
rect 571 348 572 350
rect 574 348 575 350
rect 571 343 575 348
rect 563 339 575 343
rect 563 335 567 339
rect 578 336 579 343
rect 597 366 599 368
rect 601 367 603 368
rect 638 374 644 379
rect 660 379 662 381
rect 664 379 666 381
rect 638 372 640 374
rect 642 372 644 374
rect 638 371 644 372
rect 649 373 653 375
rect 649 371 650 373
rect 652 371 653 373
rect 660 374 666 379
rect 695 379 697 381
rect 699 379 701 381
rect 695 378 701 379
rect 660 372 662 374
rect 664 372 666 374
rect 660 371 666 372
rect 601 366 611 367
rect 597 363 611 366
rect 607 359 611 363
rect 607 355 615 359
rect 611 350 615 355
rect 611 348 612 350
rect 614 348 615 350
rect 611 343 615 348
rect 603 339 615 343
rect 523 334 543 335
rect 523 332 539 334
rect 541 332 543 334
rect 523 331 543 332
rect 547 334 567 335
rect 547 332 549 334
rect 551 332 567 334
rect 547 331 567 332
rect 603 335 607 339
rect 618 336 619 343
rect 587 334 607 335
rect 587 332 589 334
rect 591 332 607 334
rect 587 331 607 332
rect 649 367 653 371
rect 672 367 696 371
rect 636 366 676 367
rect 636 364 650 366
rect 652 364 676 366
rect 636 363 676 364
rect 636 352 640 363
rect 684 362 688 364
rect 692 363 698 367
rect 684 360 685 362
rect 687 360 688 362
rect 684 359 688 360
rect 684 355 691 359
rect 634 350 640 352
rect 634 348 635 350
rect 637 348 640 350
rect 634 346 640 348
rect 644 350 648 355
rect 644 348 645 350
rect 647 348 648 350
rect 644 346 648 348
rect 636 343 640 346
rect 636 339 656 343
rect 652 335 656 339
rect 687 344 691 355
rect 694 353 698 363
rect 694 351 695 353
rect 697 351 698 353
rect 694 349 698 351
rect 687 343 705 344
rect 667 341 671 343
rect 687 342 701 343
rect 667 339 668 341
rect 670 339 671 341
rect 652 334 662 335
rect 652 332 658 334
rect 660 332 662 334
rect 652 331 662 332
rect 667 334 671 339
rect 676 341 701 342
rect 703 341 705 343
rect 676 339 678 341
rect 680 340 705 341
rect 680 339 691 340
rect 676 338 691 339
rect 667 332 668 334
rect 670 333 692 334
rect 670 332 688 333
rect 667 331 688 332
rect 690 331 692 333
rect 398 330 423 331
rect 667 330 692 331
rect 697 330 701 332
rect 181 328 182 330
rect 184 328 185 330
rect 123 327 129 328
rect 123 325 125 327
rect 127 325 129 327
rect 181 325 185 328
rect 219 328 220 330
rect 222 328 223 330
rect 389 328 390 330
rect 392 328 393 330
rect 697 328 698 330
rect 700 328 701 330
rect 219 325 223 328
rect 275 327 281 328
rect 275 325 277 327
rect 279 325 281 327
rect 389 325 393 328
rect 445 327 451 328
rect 445 325 447 327
rect 449 325 451 327
rect 639 327 645 328
rect 639 325 641 327
rect 643 325 645 327
rect 697 325 701 328
rect 123 307 125 309
rect 127 307 129 309
rect 123 306 129 307
rect 181 306 185 309
rect 181 304 182 306
rect 184 304 185 306
rect 219 306 223 309
rect 275 307 277 309
rect 279 307 281 309
rect 275 306 281 307
rect 389 306 393 309
rect 445 307 447 309
rect 449 307 451 309
rect 445 306 451 307
rect 639 307 641 309
rect 643 307 645 309
rect 639 306 645 307
rect 697 306 701 309
rect 219 304 220 306
rect 222 304 223 306
rect 389 304 390 306
rect 392 304 393 306
rect 697 304 698 306
rect 700 304 701 306
rect 151 303 176 304
rect 31 302 51 303
rect 31 300 33 302
rect 35 300 51 302
rect 31 299 51 300
rect 47 295 51 299
rect 71 302 91 303
rect 71 300 73 302
rect 75 300 91 302
rect 71 299 91 300
rect 47 291 59 295
rect 62 291 63 298
rect 55 286 59 291
rect 55 284 56 286
rect 58 284 59 286
rect 55 279 59 284
rect 51 275 59 279
rect 51 271 55 275
rect 87 295 91 299
rect 87 291 99 295
rect 102 291 103 298
rect 95 286 99 291
rect 95 284 96 286
rect 98 284 99 286
rect 95 279 99 284
rect 41 268 55 271
rect 41 266 43 268
rect 45 267 55 268
rect 45 266 47 267
rect 31 262 37 263
rect 31 260 33 262
rect 35 260 37 262
rect 31 255 37 260
rect 41 261 47 266
rect 41 259 43 261
rect 45 259 47 261
rect 41 258 47 259
rect 51 262 57 263
rect 51 260 53 262
rect 55 260 57 262
rect 31 253 33 255
rect 35 253 37 255
rect 51 255 57 260
rect 91 275 99 279
rect 91 271 95 275
rect 81 268 95 271
rect 81 266 83 268
rect 85 267 95 268
rect 85 266 87 267
rect 71 262 77 263
rect 71 260 73 262
rect 75 260 77 262
rect 51 253 53 255
rect 55 253 57 255
rect 71 255 77 260
rect 81 261 87 266
rect 81 259 83 261
rect 85 259 87 261
rect 81 258 87 259
rect 91 262 97 263
rect 91 260 93 262
rect 95 260 97 262
rect 71 253 73 255
rect 75 253 77 255
rect 91 255 97 260
rect 136 302 146 303
rect 136 300 142 302
rect 144 300 146 302
rect 136 299 146 300
rect 151 302 172 303
rect 151 300 152 302
rect 154 301 172 302
rect 174 301 176 303
rect 181 302 185 304
rect 154 300 176 301
rect 136 295 140 299
rect 120 291 140 295
rect 120 288 124 291
rect 118 286 124 288
rect 118 284 119 286
rect 121 284 124 286
rect 118 282 124 284
rect 120 271 124 282
rect 128 286 132 288
rect 151 295 155 300
rect 151 293 152 295
rect 154 293 155 295
rect 151 291 155 293
rect 160 295 175 296
rect 160 293 162 295
rect 164 294 175 295
rect 164 293 189 294
rect 160 292 185 293
rect 171 291 185 292
rect 187 291 189 293
rect 171 290 189 291
rect 128 284 129 286
rect 131 284 132 286
rect 128 279 132 284
rect 171 279 175 290
rect 168 275 175 279
rect 178 283 182 285
rect 178 281 179 283
rect 181 281 182 283
rect 168 274 172 275
rect 168 272 169 274
rect 171 272 172 274
rect 120 270 160 271
rect 168 270 172 272
rect 178 271 182 281
rect 120 268 134 270
rect 136 268 160 270
rect 120 267 160 268
rect 176 267 182 271
rect 133 263 137 267
rect 156 263 180 267
rect 122 262 128 263
rect 122 260 124 262
rect 126 260 128 262
rect 91 253 93 255
rect 95 253 97 255
rect 122 255 128 260
rect 133 261 134 263
rect 136 261 137 263
rect 133 259 137 261
rect 144 262 150 263
rect 144 260 146 262
rect 148 260 150 262
rect 122 253 124 255
rect 126 253 128 255
rect 144 255 150 260
rect 219 302 223 304
rect 228 303 253 304
rect 228 301 230 303
rect 232 302 253 303
rect 232 301 250 302
rect 228 300 250 301
rect 252 300 253 302
rect 229 295 244 296
rect 229 294 240 295
rect 215 293 240 294
rect 242 293 244 295
rect 215 291 217 293
rect 219 292 244 293
rect 249 295 253 300
rect 258 302 268 303
rect 258 300 260 302
rect 262 300 268 302
rect 258 299 268 300
rect 249 293 250 295
rect 252 293 253 295
rect 219 291 233 292
rect 249 291 253 293
rect 215 290 233 291
rect 222 283 226 285
rect 222 281 223 283
rect 225 281 226 283
rect 222 271 226 281
rect 229 279 233 290
rect 264 295 268 299
rect 264 291 284 295
rect 280 288 284 291
rect 272 286 276 288
rect 272 284 273 286
rect 275 284 276 286
rect 272 279 276 284
rect 280 286 286 288
rect 280 284 283 286
rect 285 284 286 286
rect 280 282 286 284
rect 229 275 236 279
rect 232 274 236 275
rect 232 272 233 274
rect 235 272 236 274
rect 222 267 228 271
rect 232 270 236 272
rect 280 271 284 282
rect 244 270 284 271
rect 244 268 268 270
rect 270 268 284 270
rect 244 267 284 268
rect 224 263 248 267
rect 267 263 271 267
rect 313 302 333 303
rect 313 300 329 302
rect 331 300 333 302
rect 313 299 333 300
rect 301 291 302 298
rect 313 295 317 299
rect 353 302 373 303
rect 353 300 369 302
rect 371 300 373 302
rect 353 299 373 300
rect 389 302 393 304
rect 398 303 423 304
rect 667 303 692 304
rect 398 301 400 303
rect 402 302 423 303
rect 402 301 420 302
rect 398 300 420 301
rect 422 300 423 302
rect 305 291 317 295
rect 305 286 309 291
rect 305 284 306 286
rect 308 284 309 286
rect 305 279 309 284
rect 305 275 313 279
rect 309 271 313 275
rect 309 268 323 271
rect 309 267 319 268
rect 254 262 260 263
rect 254 260 256 262
rect 258 260 260 262
rect 144 253 146 255
rect 148 253 150 255
rect 179 255 185 256
rect 179 253 181 255
rect 183 253 185 255
rect 219 255 225 256
rect 219 253 221 255
rect 223 253 225 255
rect 254 255 260 260
rect 267 261 268 263
rect 270 261 271 263
rect 267 259 271 261
rect 276 262 282 263
rect 276 260 278 262
rect 280 260 282 262
rect 254 253 256 255
rect 258 253 260 255
rect 276 255 282 260
rect 317 266 319 267
rect 321 266 323 268
rect 341 291 342 298
rect 353 295 357 299
rect 345 291 357 295
rect 345 286 349 291
rect 345 284 346 286
rect 348 284 349 286
rect 345 279 349 284
rect 345 275 353 279
rect 349 271 353 275
rect 349 268 363 271
rect 349 267 359 268
rect 307 262 313 263
rect 307 260 309 262
rect 311 260 313 262
rect 276 253 278 255
rect 280 253 282 255
rect 307 255 313 260
rect 317 261 323 266
rect 357 266 359 267
rect 361 266 363 268
rect 399 295 414 296
rect 399 294 410 295
rect 385 293 410 294
rect 412 293 414 295
rect 385 291 387 293
rect 389 292 414 293
rect 419 295 423 300
rect 428 302 438 303
rect 428 300 430 302
rect 432 300 438 302
rect 428 299 438 300
rect 419 293 420 295
rect 422 293 423 295
rect 389 291 403 292
rect 419 291 423 293
rect 385 290 403 291
rect 392 283 396 285
rect 392 281 393 283
rect 395 281 396 283
rect 392 271 396 281
rect 399 279 403 290
rect 434 295 438 299
rect 434 291 454 295
rect 450 288 454 291
rect 442 286 446 288
rect 442 284 443 286
rect 445 284 446 286
rect 442 279 446 284
rect 450 286 456 288
rect 450 284 453 286
rect 455 284 456 286
rect 450 282 456 284
rect 399 275 406 279
rect 402 274 406 275
rect 402 272 403 274
rect 405 272 406 274
rect 392 267 398 271
rect 402 270 406 272
rect 450 271 454 282
rect 414 270 454 271
rect 414 268 438 270
rect 440 268 454 270
rect 414 267 454 268
rect 317 259 319 261
rect 321 259 323 261
rect 317 258 323 259
rect 327 262 333 263
rect 327 260 329 262
rect 331 260 333 262
rect 307 253 309 255
rect 311 253 313 255
rect 327 255 333 260
rect 347 262 353 263
rect 347 260 349 262
rect 351 260 353 262
rect 327 253 329 255
rect 331 253 333 255
rect 347 255 353 260
rect 357 261 363 266
rect 394 263 418 267
rect 437 263 441 267
rect 483 302 503 303
rect 483 300 499 302
rect 501 300 503 302
rect 483 299 503 300
rect 471 291 472 298
rect 483 295 487 299
rect 523 302 543 303
rect 523 300 539 302
rect 541 300 543 302
rect 523 299 543 300
rect 547 302 567 303
rect 547 300 549 302
rect 551 300 567 302
rect 547 299 567 300
rect 475 291 487 295
rect 475 286 479 291
rect 475 284 476 286
rect 478 284 479 286
rect 475 279 479 284
rect 511 291 512 298
rect 523 295 527 299
rect 515 291 527 295
rect 475 275 483 279
rect 479 271 483 275
rect 479 268 493 271
rect 479 267 489 268
rect 357 259 359 261
rect 361 259 363 261
rect 357 258 363 259
rect 367 262 373 263
rect 367 260 369 262
rect 371 260 373 262
rect 347 253 349 255
rect 351 253 353 255
rect 367 255 373 260
rect 424 262 430 263
rect 424 260 426 262
rect 428 260 430 262
rect 367 253 369 255
rect 371 253 373 255
rect 389 255 395 256
rect 389 253 391 255
rect 393 253 395 255
rect 424 255 430 260
rect 437 261 438 263
rect 440 261 441 263
rect 437 259 441 261
rect 446 262 452 263
rect 446 260 448 262
rect 450 260 452 262
rect 424 253 426 255
rect 428 253 430 255
rect 446 255 452 260
rect 487 266 489 267
rect 491 266 493 268
rect 515 286 519 291
rect 515 284 516 286
rect 518 284 519 286
rect 515 279 519 284
rect 563 295 567 299
rect 587 302 607 303
rect 587 300 589 302
rect 591 300 607 302
rect 587 299 607 300
rect 563 291 575 295
rect 578 291 579 298
rect 571 286 575 291
rect 571 284 572 286
rect 574 284 575 286
rect 571 279 575 284
rect 515 275 523 279
rect 519 271 523 275
rect 519 268 533 271
rect 519 267 529 268
rect 477 262 483 263
rect 477 260 479 262
rect 481 260 483 262
rect 446 253 448 255
rect 450 253 452 255
rect 477 255 483 260
rect 487 261 493 266
rect 487 259 489 261
rect 491 259 493 261
rect 487 258 493 259
rect 497 262 503 263
rect 497 260 499 262
rect 501 260 503 262
rect 477 253 479 255
rect 481 253 483 255
rect 497 255 503 260
rect 527 266 529 267
rect 531 266 533 268
rect 567 275 575 279
rect 567 271 571 275
rect 603 295 607 299
rect 603 291 615 295
rect 618 291 619 298
rect 611 286 615 291
rect 611 284 612 286
rect 614 284 615 286
rect 611 279 615 284
rect 557 268 571 271
rect 557 266 559 268
rect 561 267 571 268
rect 561 266 563 267
rect 517 262 523 263
rect 517 260 519 262
rect 521 260 523 262
rect 497 253 499 255
rect 501 253 503 255
rect 517 255 523 260
rect 527 261 533 266
rect 527 259 529 261
rect 531 259 533 261
rect 527 258 533 259
rect 537 262 543 263
rect 537 260 539 262
rect 541 260 543 262
rect 517 253 519 255
rect 521 253 523 255
rect 537 255 543 260
rect 537 253 539 255
rect 541 253 543 255
rect 547 262 553 263
rect 547 260 549 262
rect 551 260 553 262
rect 547 255 553 260
rect 557 261 563 266
rect 557 259 559 261
rect 561 259 563 261
rect 557 258 563 259
rect 567 262 573 263
rect 567 260 569 262
rect 571 260 573 262
rect 547 253 549 255
rect 551 253 553 255
rect 567 255 573 260
rect 607 275 615 279
rect 607 271 611 275
rect 597 268 611 271
rect 597 266 599 268
rect 601 267 611 268
rect 601 266 603 267
rect 587 262 593 263
rect 587 260 589 262
rect 591 260 593 262
rect 567 253 569 255
rect 571 253 573 255
rect 587 255 593 260
rect 597 261 603 266
rect 597 259 599 261
rect 601 259 603 261
rect 597 258 603 259
rect 607 262 613 263
rect 607 260 609 262
rect 611 260 613 262
rect 587 253 589 255
rect 591 253 593 255
rect 607 255 613 260
rect 652 302 662 303
rect 652 300 658 302
rect 660 300 662 302
rect 652 299 662 300
rect 667 302 688 303
rect 667 300 668 302
rect 670 301 688 302
rect 690 301 692 303
rect 697 302 701 304
rect 670 300 692 301
rect 652 295 656 299
rect 636 291 656 295
rect 636 288 640 291
rect 634 286 640 288
rect 634 284 635 286
rect 637 284 640 286
rect 634 282 640 284
rect 636 271 640 282
rect 644 286 648 288
rect 667 295 671 300
rect 667 293 668 295
rect 670 293 671 295
rect 667 291 671 293
rect 676 295 691 296
rect 676 293 678 295
rect 680 294 691 295
rect 680 293 705 294
rect 676 292 701 293
rect 687 291 701 292
rect 703 291 705 293
rect 687 290 705 291
rect 644 284 645 286
rect 647 284 648 286
rect 644 279 648 284
rect 687 279 691 290
rect 684 275 691 279
rect 694 283 698 285
rect 694 281 695 283
rect 697 281 698 283
rect 684 274 688 275
rect 684 272 685 274
rect 687 272 688 274
rect 636 270 676 271
rect 684 270 688 272
rect 694 271 698 281
rect 636 268 650 270
rect 652 268 676 270
rect 636 267 676 268
rect 692 267 698 271
rect 649 263 653 267
rect 672 263 696 267
rect 638 262 644 263
rect 638 260 640 262
rect 642 260 644 262
rect 607 253 609 255
rect 611 253 613 255
rect 638 255 644 260
rect 649 261 650 263
rect 652 261 653 263
rect 649 259 653 261
rect 660 262 666 263
rect 660 260 662 262
rect 664 260 666 262
rect 638 253 640 255
rect 642 253 644 255
rect 660 255 666 260
rect 660 253 662 255
rect 664 253 666 255
rect 695 255 701 256
rect 695 253 697 255
rect 699 253 701 255
rect 82 235 84 237
rect 86 235 88 237
rect 47 231 67 232
rect 47 229 63 231
rect 65 229 67 231
rect 47 228 67 229
rect 82 230 88 235
rect 104 235 106 237
rect 108 235 110 237
rect 82 228 84 230
rect 86 228 88 230
rect 35 220 36 226
rect 47 223 51 228
rect 82 227 88 228
rect 93 229 97 231
rect 93 227 94 229
rect 96 227 97 229
rect 104 230 110 235
rect 139 235 141 237
rect 143 235 145 237
rect 139 234 145 235
rect 183 235 185 237
rect 187 235 189 237
rect 104 228 106 230
rect 108 228 110 230
rect 104 227 110 228
rect 183 230 189 235
rect 205 235 207 237
rect 209 235 211 237
rect 183 228 185 230
rect 187 228 189 230
rect 183 227 189 228
rect 194 229 198 231
rect 194 227 195 229
rect 197 227 198 229
rect 205 230 211 235
rect 240 235 242 237
rect 244 235 246 237
rect 240 234 246 235
rect 285 235 287 237
rect 289 235 291 237
rect 205 228 207 230
rect 209 228 211 230
rect 205 227 211 228
rect 285 230 291 235
rect 307 235 309 237
rect 311 235 313 237
rect 285 228 287 230
rect 289 228 291 230
rect 285 227 291 228
rect 296 229 300 231
rect 296 227 297 229
rect 299 227 300 229
rect 307 230 313 235
rect 342 235 344 237
rect 346 235 348 237
rect 342 234 348 235
rect 438 235 440 237
rect 442 235 444 237
rect 307 228 309 230
rect 311 228 313 230
rect 307 227 313 228
rect 39 219 51 223
rect 93 223 97 227
rect 116 223 140 227
rect 39 206 43 219
rect 39 204 40 206
rect 42 204 43 206
rect 39 198 43 204
rect 62 202 63 218
rect 80 222 120 223
rect 80 220 94 222
rect 96 220 120 222
rect 80 219 120 220
rect 39 194 56 198
rect 52 192 56 194
rect 41 190 47 191
rect 41 188 43 190
rect 45 188 47 190
rect 52 190 53 192
rect 55 190 56 192
rect 52 188 56 190
rect 61 192 67 193
rect 61 190 63 192
rect 65 190 67 192
rect 41 181 47 188
rect 61 181 67 190
rect 80 208 84 219
rect 128 218 132 220
rect 136 219 142 223
rect 128 216 129 218
rect 131 216 132 218
rect 128 215 132 216
rect 128 211 135 215
rect 78 206 84 208
rect 78 204 79 206
rect 81 204 84 206
rect 78 202 84 204
rect 88 206 92 211
rect 88 204 89 206
rect 91 204 92 206
rect 88 202 92 204
rect 80 199 84 202
rect 80 195 100 199
rect 96 191 100 195
rect 131 200 135 211
rect 138 209 142 219
rect 138 207 139 209
rect 141 207 142 209
rect 138 205 142 207
rect 131 199 149 200
rect 111 197 115 199
rect 131 198 145 199
rect 111 195 112 197
rect 114 195 115 197
rect 96 190 106 191
rect 96 188 102 190
rect 104 188 106 190
rect 96 187 106 188
rect 111 190 115 195
rect 120 197 145 198
rect 147 197 149 199
rect 120 195 122 197
rect 124 196 149 197
rect 124 195 135 196
rect 120 194 135 195
rect 111 188 112 190
rect 114 189 136 190
rect 114 188 132 189
rect 111 187 132 188
rect 134 187 136 189
rect 111 186 136 187
rect 141 186 145 188
rect 194 223 198 227
rect 217 223 241 227
rect 181 222 221 223
rect 181 220 195 222
rect 197 220 221 222
rect 181 219 221 220
rect 181 208 185 219
rect 229 218 233 220
rect 237 219 243 223
rect 229 216 230 218
rect 232 216 233 218
rect 229 215 233 216
rect 229 211 236 215
rect 179 206 185 208
rect 179 204 180 206
rect 182 204 185 206
rect 179 202 185 204
rect 189 206 193 211
rect 189 204 190 206
rect 192 204 193 206
rect 189 202 193 204
rect 181 199 185 202
rect 181 195 201 199
rect 197 191 201 195
rect 232 200 236 211
rect 239 209 243 219
rect 239 207 240 209
rect 242 207 243 209
rect 239 205 243 207
rect 232 199 250 200
rect 212 197 216 199
rect 232 198 246 199
rect 212 195 213 197
rect 215 195 216 197
rect 197 190 207 191
rect 197 188 203 190
rect 205 188 207 190
rect 197 187 207 188
rect 212 190 216 195
rect 221 197 246 198
rect 248 197 250 199
rect 221 195 223 197
rect 225 196 250 197
rect 225 195 236 196
rect 221 194 236 195
rect 212 188 213 190
rect 215 189 237 190
rect 215 188 233 189
rect 212 187 233 188
rect 235 187 237 189
rect 212 186 237 187
rect 242 186 246 188
rect 296 223 300 227
rect 319 223 343 227
rect 283 222 323 223
rect 283 220 297 222
rect 299 220 323 222
rect 283 219 323 220
rect 283 208 287 219
rect 331 218 335 220
rect 339 219 345 223
rect 331 216 332 218
rect 334 216 335 218
rect 331 215 335 216
rect 331 211 338 215
rect 281 206 287 208
rect 281 204 282 206
rect 284 204 287 206
rect 281 202 287 204
rect 291 206 295 211
rect 291 204 292 206
rect 294 204 295 206
rect 291 202 295 204
rect 283 199 287 202
rect 283 195 303 199
rect 299 191 303 195
rect 334 200 338 211
rect 341 209 345 219
rect 341 207 342 209
rect 344 207 345 209
rect 341 205 345 207
rect 334 199 352 200
rect 314 197 318 199
rect 334 198 348 199
rect 314 195 315 197
rect 317 195 318 197
rect 299 190 309 191
rect 299 188 305 190
rect 307 188 309 190
rect 299 187 309 188
rect 314 190 318 195
rect 323 197 348 198
rect 350 197 352 199
rect 323 195 325 197
rect 327 196 352 197
rect 327 195 338 196
rect 323 194 338 195
rect 314 188 315 190
rect 317 189 339 190
rect 317 188 335 189
rect 314 187 335 188
rect 337 187 339 189
rect 314 186 339 187
rect 344 186 348 188
rect 391 231 411 232
rect 391 229 407 231
rect 409 229 411 231
rect 391 228 411 229
rect 438 230 444 235
rect 460 235 462 237
rect 464 235 466 237
rect 438 228 440 230
rect 442 228 444 230
rect 379 220 380 226
rect 391 223 395 228
rect 438 227 444 228
rect 449 229 453 231
rect 449 227 450 229
rect 452 227 453 229
rect 460 230 466 235
rect 495 235 497 237
rect 499 235 501 237
rect 495 234 501 235
rect 539 235 541 237
rect 543 235 545 237
rect 460 228 462 230
rect 464 228 466 230
rect 460 227 466 228
rect 539 230 545 235
rect 561 235 563 237
rect 565 235 567 237
rect 539 228 541 230
rect 543 228 545 230
rect 539 227 545 228
rect 550 229 554 231
rect 550 227 551 229
rect 553 227 554 229
rect 561 230 567 235
rect 596 235 598 237
rect 600 235 602 237
rect 596 234 602 235
rect 638 235 640 237
rect 642 235 644 237
rect 561 228 563 230
rect 565 228 567 230
rect 561 227 567 228
rect 638 230 644 235
rect 660 235 662 237
rect 664 235 666 237
rect 638 228 640 230
rect 642 228 644 230
rect 638 227 644 228
rect 649 229 653 231
rect 649 227 650 229
rect 652 227 653 229
rect 660 230 666 235
rect 695 235 697 237
rect 699 235 701 237
rect 695 234 701 235
rect 660 228 662 230
rect 664 228 666 230
rect 660 227 666 228
rect 383 219 395 223
rect 449 223 453 227
rect 472 223 496 227
rect 383 206 387 219
rect 383 204 384 206
rect 386 204 387 206
rect 383 198 387 204
rect 406 202 407 218
rect 436 222 476 223
rect 436 220 450 222
rect 452 220 476 222
rect 436 219 476 220
rect 383 194 400 198
rect 396 192 400 194
rect 385 190 391 191
rect 385 188 387 190
rect 389 188 391 190
rect 396 190 397 192
rect 399 190 400 192
rect 396 188 400 190
rect 405 192 411 193
rect 405 190 407 192
rect 409 190 411 192
rect 141 184 142 186
rect 144 184 145 186
rect 242 184 243 186
rect 245 184 246 186
rect 344 184 345 186
rect 347 184 348 186
rect 83 183 89 184
rect 83 181 85 183
rect 87 181 89 183
rect 141 181 145 184
rect 184 183 190 184
rect 184 181 186 183
rect 188 181 190 183
rect 242 181 246 184
rect 286 183 292 184
rect 286 181 288 183
rect 290 181 292 183
rect 344 181 348 184
rect 385 181 391 188
rect 405 181 411 190
rect 436 208 440 219
rect 484 218 488 220
rect 492 219 498 223
rect 484 216 485 218
rect 487 216 488 218
rect 484 215 488 216
rect 484 211 491 215
rect 434 206 440 208
rect 434 204 435 206
rect 437 204 440 206
rect 434 202 440 204
rect 444 206 448 211
rect 444 204 445 206
rect 447 204 448 206
rect 444 202 448 204
rect 436 199 440 202
rect 436 195 456 199
rect 452 191 456 195
rect 487 200 491 211
rect 494 209 498 219
rect 494 207 495 209
rect 497 207 498 209
rect 494 205 498 207
rect 487 199 505 200
rect 467 197 471 199
rect 487 198 501 199
rect 467 195 468 197
rect 470 195 471 197
rect 452 190 462 191
rect 452 188 458 190
rect 460 188 462 190
rect 452 187 462 188
rect 467 190 471 195
rect 476 197 501 198
rect 503 197 505 199
rect 476 195 478 197
rect 480 196 505 197
rect 480 195 491 196
rect 476 194 491 195
rect 467 188 468 190
rect 470 189 492 190
rect 470 188 488 189
rect 467 187 488 188
rect 490 187 492 189
rect 467 186 492 187
rect 497 186 501 188
rect 550 223 554 227
rect 573 223 597 227
rect 537 222 577 223
rect 537 220 551 222
rect 553 220 577 222
rect 537 219 577 220
rect 537 208 541 219
rect 585 218 589 220
rect 593 219 599 223
rect 585 216 586 218
rect 588 216 589 218
rect 585 215 589 216
rect 585 211 592 215
rect 535 206 541 208
rect 535 204 536 206
rect 538 204 541 206
rect 535 202 541 204
rect 545 206 549 211
rect 545 204 546 206
rect 548 204 549 206
rect 545 202 549 204
rect 537 199 541 202
rect 537 195 557 199
rect 553 191 557 195
rect 588 200 592 211
rect 595 209 599 219
rect 595 207 596 209
rect 598 207 599 209
rect 595 205 599 207
rect 588 199 606 200
rect 568 197 572 199
rect 588 198 602 199
rect 568 195 569 197
rect 571 195 572 197
rect 553 190 563 191
rect 553 188 559 190
rect 561 188 563 190
rect 553 187 563 188
rect 568 190 572 195
rect 577 197 602 198
rect 604 197 606 199
rect 577 195 579 197
rect 581 196 606 197
rect 581 195 592 196
rect 577 194 592 195
rect 568 188 569 190
rect 571 189 593 190
rect 571 188 589 189
rect 568 187 589 188
rect 591 187 593 189
rect 568 186 593 187
rect 598 186 602 188
rect 649 223 653 227
rect 672 223 696 227
rect 636 222 676 223
rect 636 220 650 222
rect 652 220 676 222
rect 636 219 676 220
rect 636 208 640 219
rect 684 218 688 220
rect 692 219 698 223
rect 684 216 685 218
rect 687 216 688 218
rect 684 215 688 216
rect 684 211 691 215
rect 634 206 640 208
rect 634 204 635 206
rect 637 204 640 206
rect 634 202 640 204
rect 644 206 648 211
rect 644 204 645 206
rect 647 204 648 206
rect 644 202 648 204
rect 636 199 640 202
rect 636 195 656 199
rect 652 191 656 195
rect 687 200 691 211
rect 694 209 698 219
rect 694 207 695 209
rect 697 207 698 209
rect 694 205 698 207
rect 687 199 705 200
rect 667 197 671 199
rect 687 198 701 199
rect 667 195 668 197
rect 670 195 671 197
rect 652 190 662 191
rect 652 188 658 190
rect 660 188 662 190
rect 652 187 662 188
rect 667 190 671 195
rect 676 197 701 198
rect 703 197 705 199
rect 676 195 678 197
rect 680 196 705 197
rect 680 195 691 196
rect 676 194 691 195
rect 667 188 668 190
rect 670 189 692 190
rect 670 188 688 189
rect 667 187 688 188
rect 690 187 692 189
rect 667 186 692 187
rect 697 186 701 188
rect 497 184 498 186
rect 500 184 501 186
rect 598 184 599 186
rect 601 184 602 186
rect 697 184 698 186
rect 700 184 701 186
rect 439 183 445 184
rect 439 181 441 183
rect 443 181 445 183
rect 497 181 501 184
rect 540 183 546 184
rect 540 181 542 183
rect 544 181 546 183
rect 598 181 602 184
rect 639 183 645 184
rect 639 181 641 183
rect 643 181 645 183
rect 697 181 701 184
rect 44 163 46 165
rect 48 163 50 165
rect 44 162 50 163
rect 102 162 106 165
rect 102 160 103 162
rect 105 160 106 162
rect 72 159 97 160
rect 57 158 67 159
rect 57 156 63 158
rect 65 156 67 158
rect 57 155 67 156
rect 72 158 93 159
rect 72 156 73 158
rect 75 157 93 158
rect 95 157 97 159
rect 102 158 106 160
rect 75 156 97 157
rect 57 151 61 155
rect 41 147 61 151
rect 41 144 45 147
rect 39 142 45 144
rect 39 140 40 142
rect 42 140 45 142
rect 39 138 45 140
rect 41 127 45 138
rect 49 142 53 144
rect 72 151 76 156
rect 72 149 73 151
rect 75 149 76 151
rect 72 147 76 149
rect 81 151 96 152
rect 81 149 83 151
rect 85 150 96 151
rect 85 149 110 150
rect 81 148 106 149
rect 92 147 106 148
rect 108 147 110 149
rect 92 146 110 147
rect 49 140 50 142
rect 52 140 53 142
rect 49 135 53 140
rect 92 135 96 146
rect 89 131 96 135
rect 99 139 103 141
rect 99 137 100 139
rect 102 137 103 139
rect 89 130 93 131
rect 89 128 90 130
rect 92 128 93 130
rect 41 126 81 127
rect 89 126 93 128
rect 99 127 103 137
rect 41 124 55 126
rect 57 124 81 126
rect 41 123 81 124
rect 97 123 103 127
rect 54 119 58 123
rect 77 119 101 123
rect 43 118 49 119
rect 43 116 45 118
rect 47 116 49 118
rect 43 111 49 116
rect 54 117 55 119
rect 57 117 58 119
rect 54 115 58 117
rect 65 118 71 119
rect 65 116 67 118
rect 69 116 71 118
rect 43 109 45 111
rect 47 109 49 111
rect 65 111 71 116
rect 131 158 137 165
rect 131 156 133 158
rect 135 156 137 158
rect 131 155 137 156
rect 142 156 146 158
rect 142 154 143 156
rect 145 154 146 156
rect 142 152 146 154
rect 151 156 157 165
rect 185 163 187 165
rect 189 163 191 165
rect 185 162 191 163
rect 243 162 247 165
rect 243 160 244 162
rect 246 160 247 162
rect 285 162 289 165
rect 341 163 343 165
rect 345 163 347 165
rect 341 162 347 163
rect 285 160 286 162
rect 288 160 289 162
rect 213 159 238 160
rect 151 154 153 156
rect 155 154 157 156
rect 151 153 157 154
rect 198 158 208 159
rect 198 156 204 158
rect 206 156 208 158
rect 198 155 208 156
rect 213 158 234 159
rect 213 156 214 158
rect 216 157 234 158
rect 236 157 238 159
rect 243 158 247 160
rect 216 156 238 157
rect 129 148 146 152
rect 129 142 133 148
rect 198 151 202 155
rect 182 147 202 151
rect 182 144 186 147
rect 129 140 130 142
rect 132 140 133 142
rect 129 127 133 140
rect 152 128 153 144
rect 125 120 126 126
rect 129 123 141 127
rect 137 118 141 123
rect 180 142 186 144
rect 180 140 181 142
rect 183 140 186 142
rect 180 138 186 140
rect 182 127 186 138
rect 190 142 194 144
rect 213 151 217 156
rect 213 149 214 151
rect 216 149 217 151
rect 213 147 217 149
rect 222 151 237 152
rect 222 149 224 151
rect 226 150 237 151
rect 226 149 251 150
rect 222 148 247 149
rect 233 147 247 148
rect 249 147 251 149
rect 233 146 251 147
rect 190 140 191 142
rect 193 140 194 142
rect 190 135 194 140
rect 233 135 237 146
rect 230 131 237 135
rect 240 139 244 141
rect 240 137 241 139
rect 243 137 244 139
rect 230 130 234 131
rect 230 128 231 130
rect 233 128 234 130
rect 182 126 222 127
rect 230 126 234 128
rect 240 127 244 137
rect 182 124 196 126
rect 198 124 222 126
rect 182 123 222 124
rect 238 123 244 127
rect 195 119 199 123
rect 218 119 242 123
rect 184 118 190 119
rect 137 117 157 118
rect 137 115 153 117
rect 155 115 157 117
rect 137 114 157 115
rect 184 116 186 118
rect 188 116 190 118
rect 65 109 67 111
rect 69 109 71 111
rect 100 111 106 112
rect 100 109 102 111
rect 104 109 106 111
rect 184 111 190 116
rect 195 117 196 119
rect 198 117 199 119
rect 195 115 199 117
rect 206 118 212 119
rect 206 116 208 118
rect 210 116 212 118
rect 184 109 186 111
rect 188 109 190 111
rect 206 111 212 116
rect 285 158 289 160
rect 294 159 319 160
rect 294 157 296 159
rect 298 158 319 159
rect 298 157 316 158
rect 294 156 316 157
rect 318 156 319 158
rect 295 151 310 152
rect 295 150 306 151
rect 281 149 306 150
rect 308 149 310 151
rect 281 147 283 149
rect 285 148 310 149
rect 315 151 319 156
rect 324 158 334 159
rect 324 156 326 158
rect 328 156 334 158
rect 324 155 334 156
rect 315 149 316 151
rect 318 149 319 151
rect 285 147 299 148
rect 315 147 319 149
rect 281 146 299 147
rect 288 139 292 141
rect 288 137 289 139
rect 291 137 292 139
rect 288 127 292 137
rect 295 135 299 146
rect 330 151 334 155
rect 330 147 350 151
rect 346 144 350 147
rect 338 142 342 144
rect 338 140 339 142
rect 341 140 342 142
rect 338 135 342 140
rect 346 142 352 144
rect 346 140 349 142
rect 351 140 352 142
rect 346 138 352 140
rect 295 131 302 135
rect 298 130 302 131
rect 298 128 299 130
rect 301 128 302 130
rect 288 123 294 127
rect 298 126 302 128
rect 346 127 350 138
rect 310 126 350 127
rect 310 124 334 126
rect 336 124 350 126
rect 310 123 350 124
rect 290 119 314 123
rect 333 119 337 123
rect 385 158 391 165
rect 385 156 387 158
rect 389 156 391 158
rect 385 155 391 156
rect 396 156 400 158
rect 396 154 397 156
rect 399 154 400 156
rect 396 152 400 154
rect 405 156 411 165
rect 439 163 441 165
rect 443 163 445 165
rect 439 162 445 163
rect 497 162 501 165
rect 540 163 542 165
rect 544 163 546 165
rect 540 162 546 163
rect 598 162 602 165
rect 639 163 641 165
rect 643 163 645 165
rect 639 162 645 163
rect 697 162 701 165
rect 497 160 498 162
rect 500 160 501 162
rect 598 160 599 162
rect 601 160 602 162
rect 697 160 698 162
rect 700 160 701 162
rect 467 159 492 160
rect 405 154 407 156
rect 409 154 411 156
rect 405 153 411 154
rect 452 158 462 159
rect 452 156 458 158
rect 460 156 462 158
rect 452 155 462 156
rect 467 158 488 159
rect 467 156 468 158
rect 470 157 488 158
rect 490 157 492 159
rect 497 158 501 160
rect 568 159 593 160
rect 470 156 492 157
rect 383 148 400 152
rect 383 142 387 148
rect 383 140 384 142
rect 386 140 387 142
rect 383 127 387 140
rect 406 128 407 144
rect 379 120 380 126
rect 383 123 395 127
rect 320 118 326 119
rect 320 116 322 118
rect 324 116 326 118
rect 206 109 208 111
rect 210 109 212 111
rect 241 111 247 112
rect 241 109 243 111
rect 245 109 247 111
rect 285 111 291 112
rect 285 109 287 111
rect 289 109 291 111
rect 320 111 326 116
rect 333 117 334 119
rect 336 117 337 119
rect 333 115 337 117
rect 342 118 348 119
rect 342 116 344 118
rect 346 116 348 118
rect 320 109 322 111
rect 324 109 326 111
rect 342 111 348 116
rect 391 118 395 123
rect 452 151 456 155
rect 436 147 456 151
rect 436 144 440 147
rect 434 142 440 144
rect 434 140 435 142
rect 437 140 440 142
rect 434 138 440 140
rect 436 127 440 138
rect 444 142 448 144
rect 467 151 471 156
rect 467 149 468 151
rect 470 149 471 151
rect 467 147 471 149
rect 476 151 491 152
rect 476 149 478 151
rect 480 150 491 151
rect 480 149 505 150
rect 476 148 501 149
rect 487 147 501 148
rect 503 147 505 149
rect 487 146 505 147
rect 444 140 445 142
rect 447 140 448 142
rect 444 135 448 140
rect 487 135 491 146
rect 484 131 491 135
rect 494 139 498 141
rect 494 137 495 139
rect 497 137 498 139
rect 484 130 488 131
rect 484 128 485 130
rect 487 128 488 130
rect 436 126 476 127
rect 484 126 488 128
rect 494 127 498 137
rect 436 124 450 126
rect 452 124 476 126
rect 436 123 476 124
rect 492 123 498 127
rect 449 119 453 123
rect 472 119 496 123
rect 553 158 563 159
rect 553 156 559 158
rect 561 156 563 158
rect 553 155 563 156
rect 568 158 589 159
rect 568 156 569 158
rect 571 157 589 158
rect 591 157 593 159
rect 598 158 602 160
rect 667 159 692 160
rect 571 156 593 157
rect 553 151 557 155
rect 537 147 557 151
rect 537 144 541 147
rect 535 142 541 144
rect 535 140 536 142
rect 538 140 541 142
rect 535 138 541 140
rect 537 127 541 138
rect 545 142 549 144
rect 568 151 572 156
rect 568 149 569 151
rect 571 149 572 151
rect 568 147 572 149
rect 577 151 592 152
rect 577 149 579 151
rect 581 150 592 151
rect 581 149 606 150
rect 577 148 602 149
rect 588 147 602 148
rect 604 147 606 149
rect 588 146 606 147
rect 545 140 546 142
rect 548 140 549 142
rect 545 135 549 140
rect 588 135 592 146
rect 585 131 592 135
rect 595 139 599 141
rect 595 137 596 139
rect 598 137 599 139
rect 585 130 589 131
rect 585 128 586 130
rect 588 128 589 130
rect 537 126 577 127
rect 585 126 589 128
rect 595 127 599 137
rect 537 124 551 126
rect 553 124 577 126
rect 537 123 577 124
rect 593 123 599 127
rect 550 119 554 123
rect 573 119 597 123
rect 652 158 662 159
rect 652 156 658 158
rect 660 156 662 158
rect 652 155 662 156
rect 667 158 688 159
rect 667 156 668 158
rect 670 157 688 158
rect 690 157 692 159
rect 697 158 701 160
rect 670 156 692 157
rect 652 151 656 155
rect 636 147 656 151
rect 636 144 640 147
rect 634 142 640 144
rect 634 140 635 142
rect 637 140 640 142
rect 634 138 640 140
rect 636 127 640 138
rect 644 142 648 144
rect 667 151 671 156
rect 667 149 668 151
rect 670 149 671 151
rect 667 147 671 149
rect 676 151 691 152
rect 676 149 678 151
rect 680 150 691 151
rect 680 149 705 150
rect 676 148 701 149
rect 687 147 701 148
rect 703 147 705 149
rect 687 146 705 147
rect 644 140 645 142
rect 647 140 648 142
rect 644 135 648 140
rect 687 135 691 146
rect 684 131 691 135
rect 694 139 698 141
rect 694 137 695 139
rect 697 137 698 139
rect 684 130 688 131
rect 684 128 685 130
rect 687 128 688 130
rect 636 126 676 127
rect 684 126 688 128
rect 694 127 698 137
rect 636 124 650 126
rect 652 124 676 126
rect 636 123 676 124
rect 692 123 698 127
rect 649 119 653 123
rect 672 119 696 123
rect 438 118 444 119
rect 391 117 411 118
rect 391 115 407 117
rect 409 115 411 117
rect 391 114 411 115
rect 438 116 440 118
rect 442 116 444 118
rect 342 109 344 111
rect 346 109 348 111
rect 438 111 444 116
rect 449 117 450 119
rect 452 117 453 119
rect 449 115 453 117
rect 460 118 466 119
rect 460 116 462 118
rect 464 116 466 118
rect 438 109 440 111
rect 442 109 444 111
rect 460 111 466 116
rect 539 118 545 119
rect 539 116 541 118
rect 543 116 545 118
rect 460 109 462 111
rect 464 109 466 111
rect 495 111 501 112
rect 495 109 497 111
rect 499 109 501 111
rect 539 111 545 116
rect 550 117 551 119
rect 553 117 554 119
rect 550 115 554 117
rect 561 118 567 119
rect 561 116 563 118
rect 565 116 567 118
rect 539 109 541 111
rect 543 109 545 111
rect 561 111 567 116
rect 638 118 644 119
rect 638 116 640 118
rect 642 116 644 118
rect 561 109 563 111
rect 565 109 567 111
rect 596 111 602 112
rect 596 109 598 111
rect 600 109 602 111
rect 638 111 644 116
rect 649 117 650 119
rect 652 117 653 119
rect 649 115 653 117
rect 660 118 666 119
rect 660 116 662 118
rect 664 116 666 118
rect 638 109 640 111
rect 642 109 644 111
rect 660 111 666 116
rect 660 109 662 111
rect 664 109 666 111
rect 695 111 701 112
rect 695 109 697 111
rect 699 109 701 111
rect 82 91 84 93
rect 86 91 88 93
rect 47 87 67 88
rect 47 85 63 87
rect 65 85 67 87
rect 47 84 67 85
rect 82 86 88 91
rect 104 91 106 93
rect 108 91 110 93
rect 82 84 84 86
rect 86 84 88 86
rect 35 76 36 82
rect 47 79 51 84
rect 82 83 88 84
rect 93 85 97 87
rect 93 83 94 85
rect 96 83 97 85
rect 104 86 110 91
rect 139 91 141 93
rect 143 91 145 93
rect 139 90 145 91
rect 183 91 185 93
rect 187 91 189 93
rect 104 84 106 86
rect 108 84 110 86
rect 104 83 110 84
rect 183 86 189 91
rect 205 91 207 93
rect 209 91 211 93
rect 183 84 185 86
rect 187 84 189 86
rect 183 83 189 84
rect 194 85 198 87
rect 194 83 195 85
rect 197 83 198 85
rect 205 86 211 91
rect 240 91 242 93
rect 244 91 246 93
rect 240 90 246 91
rect 284 91 286 93
rect 288 91 290 93
rect 205 84 207 86
rect 209 84 211 86
rect 205 83 211 84
rect 284 86 290 91
rect 306 91 308 93
rect 310 91 312 93
rect 284 84 286 86
rect 288 84 290 86
rect 284 83 290 84
rect 295 85 299 87
rect 295 83 296 85
rect 298 83 299 85
rect 306 86 312 91
rect 341 91 343 93
rect 345 91 347 93
rect 341 90 347 91
rect 437 91 439 93
rect 441 91 443 93
rect 306 84 308 86
rect 310 84 312 86
rect 306 83 312 84
rect 39 75 51 79
rect 93 79 97 83
rect 116 79 140 83
rect 39 62 43 75
rect 39 60 40 62
rect 42 60 43 62
rect 39 54 43 60
rect 62 58 63 74
rect 80 78 120 79
rect 80 76 94 78
rect 96 76 120 78
rect 80 75 120 76
rect 39 50 56 54
rect 52 48 56 50
rect 41 46 47 47
rect 41 44 43 46
rect 45 44 47 46
rect 52 46 53 48
rect 55 46 56 48
rect 52 44 56 46
rect 61 48 67 49
rect 61 46 63 48
rect 65 46 67 48
rect 41 37 47 44
rect 61 37 67 46
rect 80 64 84 75
rect 128 74 132 76
rect 136 75 142 79
rect 128 72 129 74
rect 131 72 132 74
rect 128 71 132 72
rect 128 67 135 71
rect 78 62 84 64
rect 78 60 79 62
rect 81 60 84 62
rect 78 58 84 60
rect 88 62 92 67
rect 88 60 89 62
rect 91 60 92 62
rect 88 58 92 60
rect 80 55 84 58
rect 80 51 100 55
rect 96 47 100 51
rect 131 56 135 67
rect 138 65 142 75
rect 138 63 139 65
rect 141 63 142 65
rect 138 61 142 63
rect 131 55 149 56
rect 111 53 115 55
rect 131 54 145 55
rect 111 51 112 53
rect 114 51 115 53
rect 96 46 106 47
rect 96 44 102 46
rect 104 44 106 46
rect 96 43 106 44
rect 111 46 115 51
rect 120 53 145 54
rect 147 53 149 55
rect 120 51 122 53
rect 124 52 149 53
rect 124 51 135 52
rect 120 50 135 51
rect 111 44 112 46
rect 114 45 136 46
rect 114 44 132 45
rect 111 43 132 44
rect 134 43 136 45
rect 111 42 136 43
rect 141 42 145 44
rect 194 79 198 83
rect 217 79 241 83
rect 181 78 221 79
rect 181 76 195 78
rect 197 76 221 78
rect 181 75 221 76
rect 181 64 185 75
rect 229 74 233 76
rect 237 75 243 79
rect 229 72 230 74
rect 232 72 233 74
rect 229 71 233 72
rect 229 67 236 71
rect 179 62 185 64
rect 179 60 180 62
rect 182 60 185 62
rect 179 58 185 60
rect 189 62 193 67
rect 189 60 190 62
rect 192 60 193 62
rect 189 58 193 60
rect 181 55 185 58
rect 181 51 201 55
rect 197 47 201 51
rect 232 56 236 67
rect 239 65 243 75
rect 239 63 240 65
rect 242 63 243 65
rect 239 61 243 63
rect 232 55 250 56
rect 212 53 216 55
rect 232 54 246 55
rect 212 51 213 53
rect 215 51 216 53
rect 197 46 207 47
rect 197 44 203 46
rect 205 44 207 46
rect 197 43 207 44
rect 212 46 216 51
rect 221 53 246 54
rect 248 53 250 55
rect 221 51 223 53
rect 225 52 250 53
rect 225 51 236 52
rect 221 50 236 51
rect 212 44 213 46
rect 215 45 237 46
rect 215 44 233 45
rect 212 43 233 44
rect 235 43 237 45
rect 212 42 237 43
rect 242 42 246 44
rect 295 79 299 83
rect 318 79 342 83
rect 282 78 322 79
rect 282 76 296 78
rect 298 76 322 78
rect 282 75 322 76
rect 282 64 286 75
rect 330 74 334 76
rect 338 75 344 79
rect 330 72 331 74
rect 333 72 334 74
rect 330 71 334 72
rect 330 67 337 71
rect 280 62 286 64
rect 280 60 281 62
rect 283 60 286 62
rect 280 58 286 60
rect 290 62 294 67
rect 290 60 291 62
rect 293 60 294 62
rect 290 58 294 60
rect 282 55 286 58
rect 282 51 302 55
rect 298 47 302 51
rect 333 56 337 67
rect 340 65 344 75
rect 340 63 341 65
rect 343 63 344 65
rect 340 61 344 63
rect 333 55 351 56
rect 313 53 317 55
rect 333 54 347 55
rect 313 51 314 53
rect 316 51 317 53
rect 298 46 308 47
rect 298 44 304 46
rect 306 44 308 46
rect 298 43 308 44
rect 313 46 317 51
rect 322 53 347 54
rect 349 53 351 55
rect 322 51 324 53
rect 326 52 351 53
rect 326 51 337 52
rect 322 50 337 51
rect 313 44 314 46
rect 316 45 338 46
rect 316 44 334 45
rect 313 43 334 44
rect 336 43 338 45
rect 313 42 338 43
rect 343 42 347 44
rect 390 87 410 88
rect 390 85 406 87
rect 408 85 410 87
rect 390 84 410 85
rect 437 86 443 91
rect 459 91 461 93
rect 463 91 465 93
rect 437 84 439 86
rect 441 84 443 86
rect 378 76 379 82
rect 390 79 394 84
rect 437 83 443 84
rect 448 85 452 87
rect 448 83 449 85
rect 451 83 452 85
rect 459 86 465 91
rect 494 91 496 93
rect 498 91 500 93
rect 494 90 500 91
rect 538 91 540 93
rect 542 91 544 93
rect 459 84 461 86
rect 463 84 465 86
rect 459 83 465 84
rect 538 86 544 91
rect 560 91 562 93
rect 564 91 566 93
rect 538 84 540 86
rect 542 84 544 86
rect 538 83 544 84
rect 549 85 553 87
rect 549 83 550 85
rect 552 83 553 85
rect 560 86 566 91
rect 595 91 597 93
rect 599 91 601 93
rect 595 90 601 91
rect 637 91 639 93
rect 641 91 643 93
rect 560 84 562 86
rect 564 84 566 86
rect 560 83 566 84
rect 637 86 643 91
rect 659 91 661 93
rect 663 91 665 93
rect 637 84 639 86
rect 641 84 643 86
rect 637 83 643 84
rect 648 85 652 87
rect 648 83 649 85
rect 651 83 652 85
rect 659 86 665 91
rect 694 91 696 93
rect 698 91 700 93
rect 694 90 700 91
rect 659 84 661 86
rect 663 84 665 86
rect 659 83 665 84
rect 382 75 394 79
rect 448 79 452 83
rect 471 79 495 83
rect 382 62 386 75
rect 382 60 383 62
rect 385 60 386 62
rect 382 54 386 60
rect 405 58 406 74
rect 435 78 475 79
rect 435 76 449 78
rect 451 76 475 78
rect 435 75 475 76
rect 382 50 399 54
rect 395 48 399 50
rect 384 46 390 47
rect 384 44 386 46
rect 388 44 390 46
rect 395 46 396 48
rect 398 46 399 48
rect 395 44 399 46
rect 404 48 410 49
rect 404 46 406 48
rect 408 46 410 48
rect 141 40 142 42
rect 144 40 145 42
rect 242 40 243 42
rect 245 40 246 42
rect 343 40 344 42
rect 346 40 347 42
rect 83 39 89 40
rect 83 37 85 39
rect 87 37 89 39
rect 141 37 145 40
rect 184 39 190 40
rect 184 37 186 39
rect 188 37 190 39
rect 242 37 246 40
rect 285 39 291 40
rect 285 37 287 39
rect 289 37 291 39
rect 343 37 347 40
rect 384 37 390 44
rect 404 37 410 46
rect 435 64 439 75
rect 483 74 487 76
rect 491 75 497 79
rect 483 72 484 74
rect 486 72 487 74
rect 483 71 487 72
rect 483 67 490 71
rect 433 62 439 64
rect 433 60 434 62
rect 436 60 439 62
rect 433 58 439 60
rect 443 62 447 67
rect 443 60 444 62
rect 446 60 447 62
rect 443 58 447 60
rect 435 55 439 58
rect 435 51 455 55
rect 451 47 455 51
rect 486 56 490 67
rect 493 65 497 75
rect 493 63 494 65
rect 496 63 497 65
rect 493 61 497 63
rect 486 55 504 56
rect 466 53 470 55
rect 486 54 500 55
rect 466 51 467 53
rect 469 51 470 53
rect 451 46 461 47
rect 451 44 457 46
rect 459 44 461 46
rect 451 43 461 44
rect 466 46 470 51
rect 475 53 500 54
rect 502 53 504 55
rect 475 51 477 53
rect 479 52 504 53
rect 479 51 490 52
rect 475 50 490 51
rect 466 44 467 46
rect 469 45 491 46
rect 469 44 487 45
rect 466 43 487 44
rect 489 43 491 45
rect 466 42 491 43
rect 496 42 500 44
rect 549 79 553 83
rect 572 79 596 83
rect 536 78 576 79
rect 536 76 550 78
rect 552 76 576 78
rect 536 75 576 76
rect 536 64 540 75
rect 584 74 588 76
rect 592 75 598 79
rect 584 72 585 74
rect 587 72 588 74
rect 584 71 588 72
rect 584 67 591 71
rect 534 62 540 64
rect 534 60 535 62
rect 537 60 540 62
rect 534 58 540 60
rect 544 62 548 67
rect 544 60 545 62
rect 547 60 548 62
rect 544 58 548 60
rect 536 55 540 58
rect 536 51 556 55
rect 552 47 556 51
rect 587 56 591 67
rect 594 65 598 75
rect 594 63 595 65
rect 597 63 598 65
rect 594 61 598 63
rect 587 55 605 56
rect 567 53 571 55
rect 587 54 601 55
rect 567 51 568 53
rect 570 51 571 53
rect 552 46 562 47
rect 552 44 558 46
rect 560 44 562 46
rect 552 43 562 44
rect 567 46 571 51
rect 576 53 601 54
rect 603 53 605 55
rect 576 51 578 53
rect 580 52 605 53
rect 580 51 591 52
rect 576 50 591 51
rect 567 44 568 46
rect 570 45 592 46
rect 570 44 588 45
rect 567 43 588 44
rect 590 43 592 45
rect 567 42 592 43
rect 597 42 601 44
rect 648 79 652 83
rect 671 79 695 83
rect 635 78 675 79
rect 635 76 649 78
rect 651 76 675 78
rect 635 75 675 76
rect 635 64 639 75
rect 683 74 687 76
rect 691 75 697 79
rect 683 72 684 74
rect 686 72 687 74
rect 683 71 687 72
rect 683 67 690 71
rect 633 62 639 64
rect 633 60 634 62
rect 636 60 639 62
rect 633 58 639 60
rect 643 62 647 67
rect 643 60 644 62
rect 646 60 647 62
rect 643 58 647 60
rect 635 55 639 58
rect 635 51 655 55
rect 651 47 655 51
rect 686 56 690 67
rect 693 65 697 75
rect 693 63 694 65
rect 696 63 697 65
rect 693 61 697 63
rect 686 55 704 56
rect 666 53 670 55
rect 686 54 700 55
rect 666 51 667 53
rect 669 51 670 53
rect 651 46 661 47
rect 651 44 657 46
rect 659 44 661 46
rect 651 43 661 44
rect 666 46 670 51
rect 675 53 700 54
rect 702 53 704 55
rect 675 51 677 53
rect 679 52 704 53
rect 679 51 690 52
rect 675 50 690 51
rect 666 44 667 46
rect 669 45 691 46
rect 669 44 687 45
rect 666 43 687 44
rect 689 43 691 45
rect 666 42 691 43
rect 696 42 700 44
rect 496 40 497 42
rect 499 40 500 42
rect 597 40 598 42
rect 600 40 601 42
rect 696 40 697 42
rect 699 40 700 42
rect 438 39 444 40
rect 438 37 440 39
rect 442 37 444 39
rect 496 37 500 40
rect 539 39 545 40
rect 539 37 541 39
rect 543 37 545 39
rect 597 37 601 40
rect 638 39 644 40
rect 638 37 640 39
rect 642 37 644 39
rect 696 37 700 40
<< via1 >>
rect 363 388 365 390
rect 409 388 411 390
rect 454 388 456 390
rect 527 388 529 390
rect 28 384 30 386
rect 68 385 70 387
rect 106 384 108 386
rect 177 384 179 386
rect 242 384 244 386
rect 295 384 297 386
rect 330 384 332 386
rect 592 384 594 386
rect 713 385 715 387
rect 63 372 65 374
rect 41 356 43 358
rect 39 339 41 341
rect 72 356 74 358
rect 79 339 81 341
rect 103 331 105 333
rect 128 356 130 358
rect 145 339 147 341
rect 130 332 132 334
rect 192 332 194 334
rect 274 356 276 358
rect 257 339 259 341
rect 210 332 212 334
rect 272 332 274 334
rect 339 372 341 374
rect 330 356 332 358
rect 299 331 301 333
rect 323 339 325 341
rect 361 356 363 358
rect 363 339 365 341
rect 444 356 446 358
rect 427 339 429 341
rect 380 332 382 334
rect 442 332 444 334
rect 509 372 511 374
rect 500 356 502 358
rect 579 372 581 374
rect 469 331 471 333
rect 493 339 495 341
rect 531 356 533 358
rect 557 356 559 358
rect 533 339 535 341
rect 555 339 557 341
rect 588 356 590 358
rect 595 339 597 341
rect 619 331 621 333
rect 644 356 646 358
rect 661 339 663 341
rect 646 332 648 334
rect 28 316 30 318
rect 89 316 91 318
rect 153 316 155 318
rect 217 316 219 318
rect 280 316 282 318
rect 315 316 317 318
rect 347 316 349 318
rect 388 316 390 318
rect 419 316 421 318
rect 476 316 478 318
rect 566 316 568 318
rect 669 316 671 318
rect 713 316 715 318
rect 39 293 41 295
rect 41 276 43 278
rect 64 284 66 286
rect 79 293 81 295
rect 103 301 105 303
rect 72 276 74 278
rect 114 268 116 270
rect 136 284 138 286
rect 128 276 130 278
rect 192 265 194 267
rect 266 284 268 286
rect 274 276 276 278
rect 288 268 290 270
rect 210 265 212 267
rect 299 301 301 303
rect 323 293 325 295
rect 330 276 332 278
rect 363 293 365 295
rect 361 276 363 278
rect 339 263 341 265
rect 380 272 382 274
rect 460 292 462 294
rect 436 284 438 286
rect 444 276 446 278
rect 469 301 471 303
rect 493 293 495 295
rect 533 293 535 295
rect 508 284 510 286
rect 500 276 502 278
rect 555 293 557 295
rect 531 276 533 278
rect 557 276 559 278
rect 595 293 597 295
rect 619 301 621 303
rect 588 276 590 278
rect 630 268 632 270
rect 652 284 654 286
rect 644 276 646 278
rect 700 260 702 262
rect 28 243 30 245
rect 68 244 70 246
rect 106 244 108 246
rect 177 244 179 246
rect 242 244 244 246
rect 295 244 297 246
rect 330 243 332 245
rect 362 243 364 245
rect 409 244 411 246
rect 454 244 456 246
rect 713 245 715 247
rect 527 243 529 245
rect 592 243 594 245
rect 153 228 155 230
rect 53 203 55 205
rect 33 188 35 190
rect 122 212 124 214
rect 105 195 107 197
rect 210 212 212 214
rect 207 204 209 206
rect 175 188 177 190
rect 253 188 255 190
rect 291 212 293 214
rect 308 195 310 197
rect 355 188 357 190
rect 376 204 378 206
rect 399 203 401 205
rect 444 212 446 214
rect 462 204 464 206
rect 505 187 507 189
rect 545 212 547 214
rect 529 195 531 197
rect 610 203 612 205
rect 562 195 564 197
rect 644 212 646 214
rect 652 204 654 206
rect 628 195 630 197
rect 708 188 710 190
rect 25 172 27 174
rect 89 171 91 173
rect 153 172 155 174
rect 217 172 219 174
rect 280 172 282 174
rect 316 172 318 174
rect 347 172 349 174
rect 388 171 390 173
rect 419 171 421 173
rect 476 171 478 173
rect 566 172 568 174
rect 669 172 671 174
rect 713 172 715 174
rect 51 156 53 158
rect 113 156 115 158
rect 66 148 68 150
rect 83 132 85 134
rect 123 149 125 151
rect 207 149 209 151
rect 145 141 147 143
rect 255 148 257 150
rect 227 140 229 142
rect 338 156 340 158
rect 323 148 325 150
rect 340 132 342 134
rect 376 132 378 134
rect 399 141 401 143
rect 284 116 286 118
rect 462 140 464 142
rect 478 132 480 134
rect 529 149 531 151
rect 562 149 564 151
rect 610 141 612 143
rect 579 133 581 135
rect 628 149 630 151
rect 661 149 663 151
rect 678 132 680 134
rect 25 100 27 102
rect 69 101 71 103
rect 106 100 108 102
rect 177 100 179 102
rect 242 100 244 102
rect 295 100 297 102
rect 330 99 332 101
rect 363 100 365 102
rect 409 100 411 102
rect 454 100 456 102
rect 527 99 529 101
rect 592 99 594 101
rect 712 100 714 102
rect 55 59 57 61
rect 88 68 90 70
rect 106 60 108 62
rect 189 68 191 70
rect 173 51 175 53
rect 254 59 256 61
rect 206 51 208 53
rect 290 68 292 70
rect 274 51 276 53
rect 307 56 309 58
rect 375 56 377 58
rect 398 59 400 61
rect 443 68 445 70
rect 461 60 463 62
rect 544 68 546 70
rect 528 51 530 53
rect 609 59 611 61
rect 561 51 563 53
rect 643 68 645 70
rect 651 60 653 62
rect 627 51 629 53
rect 28 32 30 34
rect 89 32 91 34
rect 153 32 155 34
rect 217 32 219 34
rect 280 32 282 34
rect 316 32 318 34
rect 347 32 349 34
rect 388 32 390 34
rect 419 32 421 34
rect 476 32 478 34
rect 566 32 568 34
rect 669 32 671 34
rect 712 32 714 34
<< via2 >>
rect 363 388 365 390
rect 409 388 411 390
rect 454 388 456 390
rect 527 388 529 390
rect 28 384 30 386
rect 68 385 70 387
rect 106 384 108 386
rect 177 384 179 386
rect 242 384 244 386
rect 295 384 297 386
rect 330 384 332 386
rect 592 384 594 386
rect 713 385 715 387
rect 361 380 363 382
rect 557 380 559 382
rect 128 372 130 374
rect 274 372 276 374
rect 444 372 446 374
rect 644 372 646 374
rect 72 364 74 366
rect 500 364 502 366
rect 72 356 74 358
rect 128 356 130 358
rect 274 356 276 358
rect 361 356 363 358
rect 444 356 446 358
rect 500 356 502 358
rect 557 356 559 358
rect 644 356 646 358
rect 39 348 41 350
rect 363 348 365 350
rect 493 347 495 349
rect 595 347 597 349
rect 39 339 41 341
rect 79 339 81 341
rect 145 339 147 341
rect 257 339 259 341
rect 323 339 325 341
rect 363 339 365 341
rect 427 339 429 341
rect 493 339 495 341
rect 533 339 535 341
rect 555 339 557 341
rect 595 339 597 341
rect 661 339 663 341
rect 107 331 109 333
rect 130 332 132 334
rect 197 332 199 334
rect 210 332 212 334
rect 272 332 274 334
rect 295 331 297 333
rect 380 332 382 334
rect 442 332 444 334
rect 465 331 467 333
rect 623 331 625 333
rect 646 332 648 334
rect 28 316 30 318
rect 89 316 91 318
rect 153 316 155 318
rect 217 316 219 318
rect 280 316 282 318
rect 315 316 317 318
rect 347 316 349 318
rect 388 316 390 318
rect 419 316 421 318
rect 476 316 478 318
rect 566 316 568 318
rect 669 316 671 318
rect 713 316 715 318
rect 145 301 147 303
rect 257 301 259 303
rect 427 301 429 303
rect 661 301 663 303
rect 39 293 41 295
rect 79 293 81 295
rect 323 293 325 295
rect 363 293 365 295
rect 419 292 421 294
rect 493 293 495 295
rect 533 293 535 295
rect 555 293 557 295
rect 595 293 597 295
rect 60 284 62 286
rect 130 284 132 286
rect 209 284 211 286
rect 258 284 260 286
rect 272 284 274 286
rect 442 284 444 286
rect 519 284 521 286
rect 646 284 648 286
rect 68 276 70 278
rect 107 276 109 278
rect 169 276 171 278
rect 219 276 221 278
rect 295 276 297 278
rect 361 276 363 278
rect 465 276 467 278
rect 500 276 502 278
rect 557 276 559 278
rect 623 276 625 278
rect 370 272 372 274
rect 114 268 116 270
rect 219 268 221 270
rect 188 265 190 267
rect 614 268 616 270
rect 210 265 212 267
rect 339 263 341 265
rect 361 263 363 265
rect 557 263 559 265
rect 700 260 702 262
rect 68 255 70 257
rect 500 255 502 257
rect 28 243 30 245
rect 68 244 70 246
rect 106 244 108 246
rect 177 244 179 246
rect 242 244 244 246
rect 295 244 297 246
rect 330 243 332 245
rect 362 243 364 245
rect 409 244 411 246
rect 454 244 456 246
rect 527 243 529 245
rect 592 243 594 245
rect 713 245 715 247
rect 291 228 293 230
rect 339 228 341 230
rect 644 228 646 230
rect 258 220 260 222
rect 444 220 446 222
rect 519 220 521 222
rect 652 220 654 222
rect 161 212 163 214
rect 210 212 212 214
rect 291 212 293 214
rect 319 212 321 214
rect 419 212 421 214
rect 444 212 446 214
rect 545 212 547 214
rect 644 212 646 214
rect 53 203 55 205
rect 114 203 116 205
rect 122 203 124 205
rect 652 204 654 206
rect 113 195 115 197
rect 161 196 163 198
rect 265 196 267 198
rect 308 195 310 197
rect 33 188 35 190
rect 145 188 147 190
rect 207 188 209 190
rect 265 187 267 189
rect 319 187 321 189
rect 355 188 357 190
rect 505 187 507 189
rect 661 188 663 190
rect 380 179 382 181
rect 545 179 547 181
rect 25 172 27 174
rect 89 171 91 173
rect 153 172 155 174
rect 217 172 219 174
rect 280 172 282 174
rect 316 172 318 174
rect 347 172 349 174
rect 388 171 390 173
rect 419 171 421 173
rect 476 171 478 173
rect 566 172 568 174
rect 669 172 671 174
rect 713 172 715 174
rect 51 156 53 158
rect 113 156 115 158
rect 308 156 310 158
rect 207 149 209 151
rect 661 149 663 151
rect 145 141 147 143
rect 370 140 372 142
rect 169 132 171 134
rect 505 132 507 134
rect 614 133 616 135
rect 700 132 702 134
rect 284 116 286 118
rect 284 108 286 110
rect 651 108 653 110
rect 25 100 27 102
rect 69 101 71 103
rect 106 100 108 102
rect 177 100 179 102
rect 242 100 244 102
rect 295 100 297 102
rect 330 99 332 101
rect 363 100 365 102
rect 409 100 411 102
rect 454 100 456 102
rect 527 99 529 101
rect 592 99 594 101
rect 712 100 714 102
rect 355 90 357 92
rect 443 90 445 92
rect 61 84 63 86
rect 643 82 645 84
rect 188 76 190 78
rect 290 76 292 78
rect 33 68 35 70
rect 122 68 124 70
rect 290 68 292 70
rect 443 68 445 70
rect 544 68 546 70
rect 643 68 645 70
rect 651 60 653 62
rect 197 43 199 45
rect 544 43 546 45
rect 28 32 30 34
rect 89 32 91 34
rect 153 32 155 34
rect 217 32 219 34
rect 280 32 282 34
rect 316 32 318 34
rect 347 32 349 34
rect 388 32 390 34
rect 419 32 421 34
rect 476 32 478 34
rect 566 32 568 34
rect 669 32 671 34
rect 712 32 714 34
<< via3 >>
rect 363 388 365 390
rect 409 388 411 390
rect 454 388 456 390
rect 527 388 529 390
rect 28 384 30 386
rect 68 385 70 387
rect 106 384 108 386
rect 177 384 179 386
rect 242 384 244 386
rect 295 384 297 386
rect 330 384 332 386
rect 592 384 594 386
rect 713 385 715 387
rect 28 316 30 318
rect 89 316 91 318
rect 28 243 30 245
rect 153 316 155 318
rect 68 244 70 246
rect 106 244 108 246
rect 25 172 27 174
rect 25 100 27 102
rect 89 171 91 173
rect 69 101 71 103
rect 106 100 108 102
rect 153 172 155 174
rect 177 244 179 246
rect 177 100 179 102
rect 217 316 219 318
rect 242 244 244 246
rect 280 316 282 318
rect 315 316 317 318
rect 347 316 349 318
rect 295 244 297 246
rect 330 243 332 245
rect 362 243 364 245
rect 217 172 219 174
rect 280 172 282 174
rect 316 172 318 174
rect 347 172 349 174
rect 242 100 244 102
rect 295 100 297 102
rect 330 99 332 101
rect 388 316 390 318
rect 419 316 421 318
rect 409 244 411 246
rect 476 316 478 318
rect 566 316 568 318
rect 454 244 456 246
rect 669 316 671 318
rect 713 316 715 318
rect 527 243 529 245
rect 592 243 594 245
rect 388 171 390 173
rect 419 171 421 173
rect 476 171 478 173
rect 566 172 568 174
rect 669 172 671 174
rect 713 245 715 247
rect 713 172 715 174
rect 363 100 365 102
rect 409 100 411 102
rect 454 100 456 102
rect 527 99 529 101
rect 592 99 594 101
rect 712 100 714 102
rect 28 32 30 34
rect 89 32 91 34
rect 153 32 155 34
rect 217 32 219 34
rect 280 32 282 34
rect 316 32 318 34
rect 347 32 349 34
rect 388 32 390 34
rect 419 32 421 34
rect 476 32 478 34
rect 566 32 568 34
rect 669 32 671 34
rect 712 32 714 34
<< via4 >>
rect 5 411 7 413
rect 89 411 91 413
rect 5 316 7 318
rect 5 172 7 174
rect 5 32 7 34
rect 17 399 19 401
rect 68 399 70 401
rect 17 384 19 386
rect 28 384 30 386
rect 28 316 30 318
rect 17 243 19 245
rect 28 243 30 245
rect 25 172 27 174
rect 153 411 155 413
rect 17 100 19 102
rect 25 100 27 102
rect 28 32 30 34
rect 17 17 19 19
rect 68 17 70 19
rect 5 5 7 7
rect 106 399 108 401
rect 106 17 108 19
rect 217 411 219 413
rect 89 5 91 7
rect 177 399 179 401
rect 177 17 179 19
rect 280 411 282 413
rect 153 5 155 7
rect 242 399 244 401
rect 242 17 244 19
rect 316 411 318 413
rect 217 5 219 7
rect 295 399 297 401
rect 347 411 349 413
rect 295 17 297 19
rect 280 5 282 7
rect 330 399 332 401
rect 330 17 332 19
rect 388 411 390 413
rect 363 399 365 401
rect 316 5 318 7
rect 363 17 365 19
rect 419 411 421 413
rect 347 5 349 7
rect 409 399 411 401
rect 409 17 411 19
rect 476 411 478 413
rect 388 5 390 7
rect 454 399 456 401
rect 454 17 456 19
rect 566 411 568 413
rect 419 5 421 7
rect 527 399 529 401
rect 527 17 529 19
rect 669 411 671 413
rect 476 5 478 7
rect 592 399 594 401
rect 592 17 594 19
rect 735 411 737 413
rect 723 399 725 401
rect 713 385 715 387
rect 723 385 725 387
rect 713 316 715 318
rect 713 245 715 247
rect 723 245 725 247
rect 713 172 715 174
rect 712 100 714 102
rect 723 100 725 102
rect 566 5 568 7
rect 712 32 714 34
rect 723 17 725 19
rect 735 316 737 318
rect 735 172 737 174
rect 735 32 737 34
rect 669 5 671 7
rect 735 5 737 7
<< labels >>
rlabel alu1 113 284 113 284 1 p3
rlabel alu1 114 273 114 273 1 p3
rlabel alu1 186 261 186 261 1 p2
rlabel alu1 194 285 194 285 1 p2
rlabel alu1 186 373 186 373 1 p1
rlabel alu1 194 349 194 349 1 p1
rlabel alu1 150 385 150 385 4 vdd
rlabel alu1 150 321 150 321 4 vss
rlabel alu1 150 313 150 313 2 vss
rlabel alu1 81 277 81 277 1 b2
rlabel alu1 73 269 73 269 1 b2
rlabel alu1 89 349 89 349 1 a3
rlabel alu1 81 345 81 345 1 a3
rlabel alu1 81 357 81 357 1 b3
rlabel alu1 73 365 73 365 1 b3
rlabel alu1 89 313 89 313 2 vss
rlabel alu1 89 385 89 385 4 vdd
rlabel alu1 89 321 89 321 4 vss
rlabel alu1 65 281 65 281 1 p0
rlabel alu1 57 301 57 301 1 p0
rlabel alu1 33 365 33 365 1 b3
rlabel alu1 41 357 41 357 1 b3
rlabel alu1 49 349 49 349 1 a2
rlabel alu1 41 345 41 345 1 a2
rlabel alu1 33 269 33 269 1 b2
rlabel alu1 41 277 41 277 1 b2
rlabel alu1 49 285 49 285 1 a2
rlabel alu1 41 289 41 289 1 a2
rlabel alu1 49 313 49 313 2 vss
rlabel alu1 49 385 49 385 4 vdd
rlabel alu1 49 321 49 321 4 vss
rlabel alu1 80 289 80 289 1 a3
rlabel alu1 323 289 323 289 1 a3
rlabel alu1 323 345 323 345 1 a3
rlabel alu1 323 357 323 357 1 b1
rlabel alu1 331 365 331 365 1 b1
rlabel alu1 371 365 371 365 1 b1
rlabel via1 363 357 363 357 1 b1
rlabel alu1 331 269 331 269 1 b0
rlabel alu1 323 277 323 277 1 b0
rlabel via1 363 277 363 277 1 b0
rlabel alu1 371 269 371 269 1 b0
rlabel alu1 218 373 218 373 1 q1
rlabel alu1 210 349 210 349 1 q1
rlabel alu1 218 261 218 261 1 q2
rlabel alu1 210 285 210 285 1 q2
rlabel alu1 290 273 290 273 1 q3
rlabel alu1 291 284 291 284 1 q3
rlabel alu1 339 281 339 281 1 q0
rlabel alu1 347 301 347 301 1 q0
rlabel alu1 254 385 254 385 6 vdd
rlabel alu1 254 321 254 321 6 vss
rlabel alu1 254 313 254 313 8 vss
rlabel alu1 315 349 315 349 1 a3
rlabel alu1 315 313 315 313 8 vss
rlabel alu1 315 385 315 385 6 vdd
rlabel alu1 315 321 315 321 6 vss
rlabel alu1 355 349 355 349 1 a2
rlabel alu1 363 345 363 345 1 a2
rlabel alu1 355 285 355 285 1 a2
rlabel alu1 363 289 363 289 1 a2
rlabel alu1 355 313 355 313 8 vss
rlabel alu1 355 385 355 385 6 vdd
rlabel alu1 355 321 355 321 6 vss
rlabel alu1 493 289 493 289 1 a1
rlabel alu1 485 349 485 349 1 a1
rlabel alu1 493 345 493 345 1 a1
rlabel alu1 525 349 525 349 1 a0
rlabel alu1 533 345 533 345 1 a0
rlabel alu1 533 289 533 289 1 a0
rlabel alu1 525 285 525 285 1 a0
rlabel alu1 388 373 388 373 1 r1
rlabel alu1 380 349 380 349 1 r1
rlabel alu1 380 285 380 285 1 r2
rlabel alu1 388 261 388 261 1 r2
rlabel alu1 461 284 461 284 1 r3
rlabel alu1 460 273 460 273 1 r3
rlabel alu1 517 301 517 301 1 r0
rlabel alu1 509 281 509 281 1 r0
rlabel alu1 424 385 424 385 6 vdd
rlabel alu1 424 321 424 321 6 vss
rlabel alu1 424 313 424 313 8 vss
rlabel alu1 493 277 493 277 1 b2
rlabel alu1 501 269 501 269 1 b2
rlabel alu1 493 357 493 357 1 b3
rlabel alu1 501 365 501 365 1 b3
rlabel alu1 485 313 485 313 8 vss
rlabel alu1 485 385 485 385 6 vdd
rlabel alu1 485 321 485 321 6 vss
rlabel alu1 541 365 541 365 1 b3
rlabel alu1 533 357 533 357 1 b3
rlabel alu1 541 269 541 269 1 b2
rlabel alu1 533 277 533 277 1 b2
rlabel alu1 525 313 525 313 8 vss
rlabel alu1 525 385 525 385 6 vdd
rlabel alu1 525 321 525 321 6 vss
rlabel alu1 596 289 596 289 1 a1
rlabel alu1 605 349 605 349 1 a1
rlabel alu1 597 345 597 345 1 a1
rlabel alu1 597 357 597 357 1 b1
rlabel alu1 589 365 589 365 1 b1
rlabel alu1 549 365 549 365 1 b1
rlabel via1 557 357 557 357 1 b1
rlabel alu1 565 349 565 349 1 a0
rlabel alu1 557 345 557 345 1 a0
rlabel alu1 597 277 597 277 1 b0
rlabel alu1 589 269 589 269 1 b0
rlabel via1 557 277 557 277 1 b0
rlabel alu1 549 269 549 269 1 b0
rlabel alu1 557 289 557 289 1 a0
rlabel alu1 565 285 565 285 1 a0
rlabel alu1 702 373 702 373 1 o1
rlabel alu1 710 349 710 349 1 o1
rlabel alu1 702 261 702 261 1 s2
rlabel alu1 629 284 629 284 1 s3
rlabel alu1 630 273 630 273 1 s3
rlabel alu1 573 301 573 301 1 o0
rlabel alu1 581 281 581 281 1 o0
rlabel alu1 666 385 666 385 4 vdd
rlabel alu1 666 321 666 321 4 vss
rlabel alu1 666 313 666 313 2 vss
rlabel alu1 605 313 605 313 2 vss
rlabel alu1 605 385 605 385 4 vdd
rlabel alu1 605 321 605 321 4 vss
rlabel alu1 565 313 565 313 2 vss
rlabel alu1 565 385 565 385 4 vdd
rlabel alu1 565 321 565 321 4 vss
rlabel alu1 710 285 710 285 1 s2
rlabel alu1 709 64 709 64 1 o4
rlabel alu1 661 69 661 69 1 p0
rlabel alu1 661 57 661 57 1 u0
rlabel alu1 665 97 665 97 4 vdd
rlabel alu1 665 33 665 33 4 vss
rlabel alu1 666 177 666 177 4 vss
rlabel alu1 666 241 666 241 4 vdd
rlabel alu1 662 201 662 201 1 r0
rlabel alu1 654 205 654 205 1 r0
rlabel pmos 646 213 646 213 1 q0
rlabel alu1 654 213 654 213 1 q0
rlabel alu1 662 213 662 213 1 q0
rlabel alu1 670 213 670 213 1 q0
rlabel alu1 678 209 678 209 1 q0
rlabel alu1 666 169 666 169 2 vss
rlabel alu1 666 105 666 105 2 vdd
rlabel alu1 661 133 661 133 1 s2
rlabel alu1 671 133 671 133 1 s2
rlabel alu1 710 208 710 208 1 t5
rlabel alu1 629 142 629 142 1 t4
rlabel alu1 629 208 629 208 1 t3
rlabel alu1 641 189 641 189 1 t3
rlabel alu1 710 142 710 142 1 o2
rlabel alu1 565 133 565 133 1 s3
rlabel alu1 567 169 567 169 2 vss
rlabel alu1 567 105 567 105 2 vdd
rlabel pmos 547 213 547 213 1 r1
rlabel alu1 555 213 555 213 1 r1
rlabel alu1 563 213 563 213 1 r1
rlabel alu1 571 213 571 213 1 r1
rlabel alu1 579 209 579 209 1 r1
rlabel alu1 567 177 567 177 4 vss
rlabel alu1 567 241 567 241 4 vdd
rlabel alu1 566 97 566 97 4 vdd
rlabel alu1 566 33 566 33 4 vss
rlabel alu1 561 69 561 69 1 p1
rlabel alu1 510 134 510 134 1 o3
rlabel alu1 510 208 510 208 1 t6
rlabel alu1 466 169 466 169 2 vss
rlabel alu1 466 105 466 105 2 vdd
rlabel alu1 478 209 478 209 1 q1
rlabel alu1 470 213 470 213 1 q1
rlabel alu1 462 213 462 213 1 q1
rlabel alu1 454 213 454 213 1 q1
rlabel pmos 446 213 446 213 1 q1
rlabel alu1 466 177 466 177 4 vss
rlabel alu1 466 241 466 241 4 vdd
rlabel alu1 465 97 465 97 4 vdd
rlabel alu1 465 33 465 33 4 vss
rlabel alu1 462 69 462 69 1 u1
rlabel alu1 509 66 509 66 1 o5
rlabel alu1 377 136 377 136 1 t2
rlabel alu1 377 208 377 208 1 t1
rlabel alu1 393 105 393 105 8 vdd
rlabel alu1 393 169 393 169 8 vss
rlabel alu1 393 241 393 241 6 vdd
rlabel alu1 393 177 393 177 6 vss
rlabel alu1 392 33 392 33 6 vss
rlabel alu1 392 97 392 97 6 vdd
rlabel alu1 357 199 357 199 1 u1
rlabel alu1 276 134 276 134 1 u0
rlabel alu1 313 241 313 241 4 vdd
rlabel alu1 313 177 313 177 4 vss
rlabel alu1 320 105 320 105 8 vdd
rlabel alu1 320 169 320 169 8 vss
rlabel alu1 356 65 356 65 1 o6
rlabel alu1 308 69 308 69 1 p2
rlabel alu1 312 97 312 97 4 vdd
rlabel alu1 312 33 312 33 4 vss
rlabel alu1 216 133 216 133 1 r2
rlabel alu1 208 133 208 133 1 r2
rlabel alu1 200 133 200 133 1 r2
rlabel pmos 192 133 192 133 1 r2
rlabel alu1 223 209 223 209 1 q2
rlabel alu1 215 213 215 213 1 q2
rlabel alu1 207 213 207 213 1 q2
rlabel alu1 199 213 199 213 1 q2
rlabel pmos 191 213 191 213 1 q2
rlabel alu1 211 177 211 177 4 vss
rlabel alu1 211 241 211 241 4 vdd
rlabel alu1 212 105 212 105 2 vdd
rlabel alu1 212 169 212 169 2 vss
rlabel alu1 208 69 208 69 1 p3
rlabel alu1 211 33 211 33 4 vss
rlabel alu1 211 97 211 97 4 vdd
rlabel alu1 33 209 33 209 1 ca1
rlabel alu1 122 209 122 209 1 r3
rlabel alu1 114 213 114 213 1 r3
rlabel alu1 106 213 106 213 1 r3
rlabel alu1 98 213 98 213 1 r3
rlabel pmos 90 213 90 213 1 r3
rlabel alu1 75 133 75 133 1 q3
rlabel alu1 67 133 67 133 1 q3
rlabel alu1 59 133 59 133 1 q3
rlabel pmos 51 133 51 133 1 q3
rlabel alu1 139 105 139 105 8 vdd
rlabel alu1 139 169 139 169 8 vss
rlabel alu1 131 117 131 117 8 z
rlabel alu1 123 137 123 137 8 z
rlabel alu1 71 105 71 105 2 vdd
rlabel alu1 71 169 71 169 2 vss
rlabel alu0 82 209 82 209 4 con
rlabel alu1 110 177 110 177 4 vss
rlabel alu1 110 241 110 241 4 vdd
rlabel alu1 49 241 49 241 6 vdd
rlabel alu1 49 177 49 177 6 vss
rlabel alu1 154 65 154 65 1 o7
rlabel alu1 108 69 108 69 1 ca1
rlabel alu1 110 33 110 33 4 vss
rlabel alu1 110 97 110 97 4 vdd
rlabel alu1 49 97 49 97 6 vdd
rlabel alu1 49 33 49 33 6 vss
rlabel alu1 628 57 628 57 1 x1
rlabel alu1 376 66 376 66 1 x2
rlabel alu1 275 62 275 62 1 x3
rlabel alu1 33 63 33 63 1 ca3
<< end >>
