magic
tech scmos
timestamp 1508926407
<< ab >>
rect 5 -68 45 76
rect 47 -4 53 12
rect 55 -68 95 76
rect 97 -4 103 12
rect 97 -68 103 -60
rect 105 -68 201 76
<< nwell >>
rect 0 36 206 81
rect 0 -73 206 -28
<< pwell >>
rect 0 -28 206 36
<< poly >>
rect 14 70 16 74
rect 24 70 26 74
rect 34 70 36 74
rect 64 70 66 74
rect 74 70 76 74
rect 84 70 86 74
rect 122 70 124 74
rect 132 70 134 74
rect 142 70 144 74
rect 14 47 16 51
rect 10 45 16 47
rect 10 43 12 45
rect 14 43 16 45
rect 10 41 16 43
rect 14 30 16 41
rect 24 39 26 51
rect 64 47 66 51
rect 60 45 66 47
rect 60 43 62 45
rect 64 43 66 45
rect 34 39 36 42
rect 60 41 66 43
rect 20 37 26 39
rect 20 35 22 37
rect 24 35 26 37
rect 20 33 26 35
rect 30 37 36 39
rect 30 35 32 37
rect 34 35 36 37
rect 30 33 36 35
rect 21 30 23 33
rect 34 30 36 33
rect 64 30 66 41
rect 74 39 76 51
rect 160 67 162 72
rect 167 67 169 72
rect 190 70 192 74
rect 177 58 179 63
rect 177 42 179 45
rect 84 39 86 42
rect 122 39 124 42
rect 132 39 134 42
rect 142 39 144 42
rect 160 39 162 42
rect 167 39 169 42
rect 177 40 186 42
rect 70 37 76 39
rect 70 35 72 37
rect 74 35 76 37
rect 70 33 76 35
rect 80 37 86 39
rect 80 35 82 37
rect 84 35 86 37
rect 80 33 86 35
rect 120 37 126 39
rect 120 35 122 37
rect 124 35 126 37
rect 120 33 126 35
rect 130 37 136 39
rect 130 35 132 37
rect 134 35 136 37
rect 130 33 136 35
rect 140 37 162 39
rect 140 35 142 37
rect 144 35 149 37
rect 151 35 162 37
rect 140 33 162 35
rect 166 37 172 39
rect 166 35 168 37
rect 170 35 172 37
rect 166 33 172 35
rect 71 30 73 33
rect 84 30 86 33
rect 14 12 16 17
rect 21 12 23 17
rect 34 11 36 16
rect 64 12 66 17
rect 71 12 73 17
rect 122 24 124 33
rect 133 30 135 33
rect 140 30 142 33
rect 160 30 162 33
rect 170 30 172 33
rect 180 38 182 40
rect 184 38 186 40
rect 180 36 186 38
rect 84 11 86 16
rect 180 23 182 36
rect 190 32 192 45
rect 186 30 192 32
rect 186 28 188 30
rect 190 28 192 30
rect 186 26 192 28
rect 190 23 192 26
rect 160 11 162 16
rect 170 11 172 16
rect 122 6 124 10
rect 133 6 135 10
rect 140 6 142 10
rect 180 8 182 13
rect 190 6 192 10
rect 122 -2 124 2
rect 133 -2 135 2
rect 140 -2 142 2
rect 14 -9 16 -4
rect 21 -9 23 -4
rect 34 -8 36 -3
rect 64 -9 66 -4
rect 71 -9 73 -4
rect 84 -8 86 -3
rect 14 -33 16 -22
rect 21 -25 23 -22
rect 34 -25 36 -22
rect 20 -27 26 -25
rect 20 -29 22 -27
rect 24 -29 26 -27
rect 20 -31 26 -29
rect 30 -27 36 -25
rect 30 -29 32 -27
rect 34 -29 36 -27
rect 30 -31 36 -29
rect 10 -35 16 -33
rect 10 -37 12 -35
rect 14 -37 16 -35
rect 10 -39 16 -37
rect 14 -43 16 -39
rect 24 -43 26 -31
rect 34 -34 36 -31
rect 64 -33 66 -22
rect 71 -25 73 -22
rect 84 -25 86 -22
rect 122 -25 124 -16
rect 160 -8 162 -3
rect 170 -8 172 -3
rect 180 -5 182 0
rect 190 -2 192 2
rect 133 -25 135 -22
rect 140 -25 142 -22
rect 160 -25 162 -22
rect 170 -25 172 -22
rect 70 -27 76 -25
rect 70 -29 72 -27
rect 74 -29 76 -27
rect 70 -31 76 -29
rect 80 -27 86 -25
rect 80 -29 82 -27
rect 84 -29 86 -27
rect 80 -31 86 -29
rect 120 -27 126 -25
rect 120 -29 122 -27
rect 124 -29 126 -27
rect 120 -31 126 -29
rect 130 -27 136 -25
rect 130 -29 132 -27
rect 134 -29 136 -27
rect 130 -31 136 -29
rect 140 -27 162 -25
rect 140 -29 142 -27
rect 144 -29 149 -27
rect 151 -29 162 -27
rect 140 -31 162 -29
rect 166 -27 172 -25
rect 166 -29 168 -27
rect 170 -29 172 -27
rect 166 -31 172 -29
rect 180 -28 182 -15
rect 190 -18 192 -15
rect 186 -20 192 -18
rect 186 -22 188 -20
rect 190 -22 192 -20
rect 186 -24 192 -22
rect 180 -30 186 -28
rect 60 -35 66 -33
rect 60 -37 62 -35
rect 64 -37 66 -35
rect 60 -39 66 -37
rect 64 -43 66 -39
rect 74 -43 76 -31
rect 84 -34 86 -31
rect 122 -34 124 -31
rect 132 -34 134 -31
rect 142 -34 144 -31
rect 160 -34 162 -31
rect 167 -34 169 -31
rect 180 -32 182 -30
rect 184 -32 186 -30
rect 177 -34 186 -32
rect 177 -37 179 -34
rect 190 -37 192 -24
rect 177 -55 179 -50
rect 14 -66 16 -62
rect 24 -66 26 -62
rect 34 -66 36 -62
rect 64 -66 66 -62
rect 74 -66 76 -62
rect 84 -66 86 -62
rect 122 -66 124 -62
rect 132 -66 134 -62
rect 142 -66 144 -62
rect 160 -64 162 -59
rect 167 -64 169 -59
rect 190 -66 192 -62
<< ndif >>
rect 9 23 14 30
rect 7 21 14 23
rect 7 19 9 21
rect 11 19 14 21
rect 7 17 14 19
rect 16 17 21 30
rect 23 17 34 30
rect 25 16 34 17
rect 36 28 43 30
rect 36 26 39 28
rect 41 26 43 28
rect 36 20 43 26
rect 59 23 64 30
rect 36 18 39 20
rect 41 18 43 20
rect 36 16 43 18
rect 57 21 64 23
rect 57 19 59 21
rect 61 19 64 21
rect 57 17 64 19
rect 66 17 71 30
rect 73 17 84 30
rect 25 11 32 16
rect 75 16 84 17
rect 86 28 93 30
rect 86 26 89 28
rect 91 26 93 28
rect 86 20 93 26
rect 126 24 133 30
rect 86 18 89 20
rect 91 18 93 20
rect 86 16 93 18
rect 115 21 122 24
rect 115 19 117 21
rect 119 19 122 21
rect 115 17 122 19
rect 75 11 82 16
rect 25 9 28 11
rect 30 9 32 11
rect 25 7 32 9
rect 75 9 78 11
rect 80 9 82 11
rect 117 10 122 17
rect 124 14 133 24
rect 124 12 128 14
rect 130 12 133 14
rect 124 10 133 12
rect 135 10 140 30
rect 142 23 147 30
rect 153 28 160 30
rect 153 26 155 28
rect 157 26 160 28
rect 142 21 149 23
rect 142 19 145 21
rect 147 19 149 21
rect 142 17 149 19
rect 153 21 160 26
rect 153 19 155 21
rect 157 19 160 21
rect 142 10 147 17
rect 153 16 160 19
rect 162 28 170 30
rect 162 26 165 28
rect 167 26 170 28
rect 162 16 170 26
rect 172 23 177 30
rect 172 20 180 23
rect 172 18 175 20
rect 177 18 180 20
rect 172 16 180 18
rect 175 13 180 16
rect 182 17 190 23
rect 182 15 185 17
rect 187 15 190 17
rect 182 13 190 15
rect 75 7 82 9
rect 185 10 190 13
rect 192 21 199 23
rect 192 19 195 21
rect 197 19 199 21
rect 192 17 199 19
rect 192 10 197 17
rect 25 -1 32 1
rect 25 -3 28 -1
rect 30 -3 32 -1
rect 75 -1 82 1
rect 75 -3 78 -1
rect 80 -3 82 -1
rect 25 -8 32 -3
rect 25 -9 34 -8
rect 7 -11 14 -9
rect 7 -13 9 -11
rect 11 -13 14 -11
rect 7 -15 14 -13
rect 9 -22 14 -15
rect 16 -22 21 -9
rect 23 -22 34 -9
rect 36 -10 43 -8
rect 75 -8 82 -3
rect 75 -9 84 -8
rect 36 -12 39 -10
rect 41 -12 43 -10
rect 36 -18 43 -12
rect 57 -11 64 -9
rect 57 -13 59 -11
rect 61 -13 64 -11
rect 57 -15 64 -13
rect 36 -20 39 -18
rect 41 -20 43 -18
rect 36 -22 43 -20
rect 59 -22 64 -15
rect 66 -22 71 -9
rect 73 -22 84 -9
rect 86 -10 93 -8
rect 117 -9 122 -2
rect 86 -12 89 -10
rect 91 -12 93 -10
rect 86 -18 93 -12
rect 115 -11 122 -9
rect 115 -13 117 -11
rect 119 -13 122 -11
rect 115 -16 122 -13
rect 124 -4 133 -2
rect 124 -6 128 -4
rect 130 -6 133 -4
rect 124 -16 133 -6
rect 86 -20 89 -18
rect 91 -20 93 -18
rect 86 -22 93 -20
rect 126 -22 133 -16
rect 135 -22 140 -2
rect 142 -9 147 -2
rect 185 -5 190 -2
rect 175 -8 180 -5
rect 142 -11 149 -9
rect 142 -13 145 -11
rect 147 -13 149 -11
rect 142 -15 149 -13
rect 153 -11 160 -8
rect 153 -13 155 -11
rect 157 -13 160 -11
rect 142 -22 147 -15
rect 153 -18 160 -13
rect 153 -20 155 -18
rect 157 -20 160 -18
rect 153 -22 160 -20
rect 162 -18 170 -8
rect 162 -20 165 -18
rect 167 -20 170 -18
rect 162 -22 170 -20
rect 172 -10 180 -8
rect 172 -12 175 -10
rect 177 -12 180 -10
rect 172 -15 180 -12
rect 182 -7 190 -5
rect 182 -9 185 -7
rect 187 -9 190 -7
rect 182 -15 190 -9
rect 192 -9 197 -2
rect 192 -11 199 -9
rect 192 -13 195 -11
rect 197 -13 199 -11
rect 192 -15 199 -13
rect 172 -22 177 -15
<< pdif >>
rect 7 68 14 70
rect 7 66 9 68
rect 11 66 14 68
rect 7 61 14 66
rect 7 59 9 61
rect 11 59 14 61
rect 7 51 14 59
rect 16 62 24 70
rect 16 60 19 62
rect 21 60 24 62
rect 16 55 24 60
rect 16 53 19 55
rect 21 53 24 55
rect 16 51 24 53
rect 26 68 34 70
rect 26 66 29 68
rect 31 66 34 68
rect 26 61 34 66
rect 26 59 29 61
rect 31 59 34 61
rect 26 51 34 59
rect 28 42 34 51
rect 36 63 41 70
rect 57 68 64 70
rect 57 66 59 68
rect 61 66 64 68
rect 36 61 43 63
rect 36 59 39 61
rect 41 59 43 61
rect 36 54 43 59
rect 36 52 39 54
rect 41 52 43 54
rect 36 50 43 52
rect 57 61 64 66
rect 57 59 59 61
rect 61 59 64 61
rect 57 51 64 59
rect 66 62 74 70
rect 66 60 69 62
rect 71 60 74 62
rect 66 55 74 60
rect 66 53 69 55
rect 71 53 74 55
rect 66 51 74 53
rect 76 68 84 70
rect 76 66 79 68
rect 81 66 84 68
rect 76 61 84 66
rect 76 59 79 61
rect 81 59 84 61
rect 76 51 84 59
rect 36 42 41 50
rect 78 42 84 51
rect 86 63 91 70
rect 86 61 93 63
rect 86 59 89 61
rect 91 59 93 61
rect 86 54 93 59
rect 117 55 122 70
rect 86 52 89 54
rect 91 52 93 54
rect 86 50 93 52
rect 115 53 122 55
rect 115 51 117 53
rect 119 51 122 53
rect 86 42 91 50
rect 115 46 122 51
rect 115 44 117 46
rect 119 44 122 46
rect 115 42 122 44
rect 124 68 132 70
rect 124 66 127 68
rect 129 66 132 68
rect 124 61 132 66
rect 124 59 127 61
rect 129 59 132 61
rect 124 42 132 59
rect 134 60 142 70
rect 134 58 137 60
rect 139 58 142 60
rect 134 53 142 58
rect 134 51 137 53
rect 139 51 142 53
rect 134 42 142 51
rect 144 68 158 70
rect 144 66 149 68
rect 151 67 158 68
rect 181 68 190 70
rect 151 66 160 67
rect 144 61 160 66
rect 144 59 149 61
rect 151 59 160 61
rect 144 42 160 59
rect 162 42 167 67
rect 169 58 174 67
rect 181 66 184 68
rect 186 66 190 68
rect 181 58 190 66
rect 169 49 177 58
rect 169 47 172 49
rect 174 47 177 49
rect 169 45 177 47
rect 179 45 190 58
rect 192 58 197 70
rect 192 56 199 58
rect 192 54 195 56
rect 197 54 199 56
rect 192 49 199 54
rect 192 47 195 49
rect 197 47 199 49
rect 192 45 199 47
rect 169 42 174 45
rect 28 -43 34 -34
rect 7 -51 14 -43
rect 7 -53 9 -51
rect 11 -53 14 -51
rect 7 -58 14 -53
rect 7 -60 9 -58
rect 11 -60 14 -58
rect 7 -62 14 -60
rect 16 -45 24 -43
rect 16 -47 19 -45
rect 21 -47 24 -45
rect 16 -52 24 -47
rect 16 -54 19 -52
rect 21 -54 24 -52
rect 16 -62 24 -54
rect 26 -51 34 -43
rect 26 -53 29 -51
rect 31 -53 34 -51
rect 26 -58 34 -53
rect 26 -60 29 -58
rect 31 -60 34 -58
rect 26 -62 34 -60
rect 36 -42 41 -34
rect 36 -44 43 -42
rect 78 -43 84 -34
rect 36 -46 39 -44
rect 41 -46 43 -44
rect 36 -51 43 -46
rect 36 -53 39 -51
rect 41 -53 43 -51
rect 36 -55 43 -53
rect 57 -51 64 -43
rect 57 -53 59 -51
rect 61 -53 64 -51
rect 36 -62 41 -55
rect 57 -58 64 -53
rect 57 -60 59 -58
rect 61 -60 64 -58
rect 57 -62 64 -60
rect 66 -45 74 -43
rect 66 -47 69 -45
rect 71 -47 74 -45
rect 66 -52 74 -47
rect 66 -54 69 -52
rect 71 -54 74 -52
rect 66 -62 74 -54
rect 76 -51 84 -43
rect 76 -53 79 -51
rect 81 -53 84 -51
rect 76 -58 84 -53
rect 76 -60 79 -58
rect 81 -60 84 -58
rect 76 -62 84 -60
rect 86 -42 91 -34
rect 115 -36 122 -34
rect 115 -38 117 -36
rect 119 -38 122 -36
rect 86 -44 93 -42
rect 86 -46 89 -44
rect 91 -46 93 -44
rect 86 -51 93 -46
rect 115 -43 122 -38
rect 115 -45 117 -43
rect 119 -45 122 -43
rect 115 -47 122 -45
rect 86 -53 89 -51
rect 91 -53 93 -51
rect 86 -55 93 -53
rect 86 -62 91 -55
rect 117 -62 122 -47
rect 124 -51 132 -34
rect 124 -53 127 -51
rect 129 -53 132 -51
rect 124 -58 132 -53
rect 124 -60 127 -58
rect 129 -60 132 -58
rect 124 -62 132 -60
rect 134 -43 142 -34
rect 134 -45 137 -43
rect 139 -45 142 -43
rect 134 -50 142 -45
rect 134 -52 137 -50
rect 139 -52 142 -50
rect 134 -62 142 -52
rect 144 -51 160 -34
rect 144 -53 149 -51
rect 151 -53 160 -51
rect 144 -58 160 -53
rect 144 -60 149 -58
rect 151 -59 160 -58
rect 162 -59 167 -34
rect 169 -37 174 -34
rect 169 -39 177 -37
rect 169 -41 172 -39
rect 174 -41 177 -39
rect 169 -50 177 -41
rect 179 -50 190 -37
rect 169 -59 174 -50
rect 181 -58 190 -50
rect 151 -60 158 -59
rect 144 -62 158 -60
rect 181 -60 184 -58
rect 186 -60 190 -58
rect 181 -62 190 -60
rect 192 -39 199 -37
rect 192 -41 195 -39
rect 197 -41 199 -39
rect 192 -46 199 -41
rect 192 -48 195 -46
rect 197 -48 199 -46
rect 192 -50 199 -48
rect 192 -62 197 -50
<< alu1 >>
rect 3 72 203 76
rect -11 68 203 72
rect -11 -60 -7 68
rect 38 61 43 63
rect 38 59 39 61
rect 41 59 43 61
rect 7 46 11 55
rect 38 54 43 59
rect 88 61 93 63
rect 88 59 89 61
rect 91 59 93 61
rect 38 52 39 54
rect 41 52 43 54
rect 38 50 43 52
rect 7 45 20 46
rect 7 43 12 45
rect 14 43 17 45
rect 19 43 20 45
rect 7 42 20 43
rect 14 37 28 38
rect 14 35 22 37
rect 24 35 28 37
rect 14 34 28 35
rect 14 28 19 34
rect 14 26 15 28
rect 17 26 19 28
rect 14 25 19 26
rect 39 28 43 50
rect 57 46 61 55
rect 88 54 93 59
rect 186 58 199 62
rect 88 52 89 54
rect 91 52 93 54
rect 88 50 93 52
rect 57 45 70 46
rect 57 43 58 45
rect 60 43 62 45
rect 64 43 70 45
rect 57 42 70 43
rect 41 26 43 28
rect 39 23 43 26
rect 64 37 78 38
rect 64 35 72 37
rect 74 35 78 37
rect 64 34 78 35
rect 64 28 69 34
rect 64 26 65 28
rect 67 26 69 28
rect 64 25 69 26
rect 31 20 43 23
rect 89 28 93 50
rect 91 26 93 28
rect 89 23 93 26
rect 31 18 39 20
rect 41 18 43 20
rect 81 20 93 23
rect 81 18 89 20
rect 91 18 93 20
rect 114 53 120 55
rect 194 56 199 58
rect 194 54 195 56
rect 197 54 199 56
rect 114 51 117 53
rect 119 51 120 53
rect 114 46 120 51
rect 114 44 117 46
rect 119 44 120 46
rect 114 42 120 44
rect 114 22 118 42
rect 130 45 168 46
rect 130 43 131 45
rect 133 43 168 45
rect 130 42 168 43
rect 163 39 168 42
rect 138 37 153 38
rect 138 35 142 37
rect 144 35 149 37
rect 151 35 153 37
rect 138 34 153 35
rect 163 37 171 39
rect 163 35 168 37
rect 170 35 171 37
rect 147 28 151 34
rect 163 33 171 35
rect 194 49 199 54
rect 194 47 195 49
rect 197 47 199 49
rect 194 45 199 47
rect 147 26 148 28
rect 150 26 151 28
rect 147 25 151 26
rect 114 21 136 22
rect 114 19 117 21
rect 119 19 133 21
rect 135 19 136 21
rect 114 18 136 19
rect 195 23 199 45
rect 194 21 199 23
rect 194 19 195 21
rect 197 19 199 21
rect 31 17 43 18
rect 81 17 93 18
rect 194 17 199 19
rect 3 11 203 12
rect 3 9 28 11
rect 30 9 78 11
rect 80 9 203 11
rect 3 -1 203 9
rect 3 -3 28 -1
rect 30 -3 78 -1
rect 80 -3 203 -1
rect 3 -4 203 -3
rect 31 -10 43 -9
rect 81 -10 93 -9
rect 14 -18 19 -17
rect 14 -20 15 -18
rect 17 -20 19 -18
rect 14 -26 19 -20
rect 31 -12 39 -10
rect 41 -12 43 -10
rect 31 -15 43 -12
rect 39 -18 43 -15
rect 41 -20 43 -18
rect 14 -27 28 -26
rect 14 -29 22 -27
rect 24 -29 28 -27
rect 14 -30 28 -29
rect 7 -35 20 -34
rect 7 -37 12 -35
rect 14 -37 17 -35
rect 19 -37 20 -35
rect 7 -38 20 -37
rect 7 -47 11 -38
rect 39 -42 43 -20
rect 64 -18 69 -17
rect 64 -20 65 -18
rect 67 -20 69 -18
rect 64 -26 69 -20
rect 81 -12 89 -10
rect 91 -12 93 -10
rect 81 -15 93 -12
rect 89 -18 93 -15
rect 91 -20 93 -18
rect 64 -27 78 -26
rect 64 -29 72 -27
rect 74 -29 78 -27
rect 64 -30 78 -29
rect 38 -44 43 -42
rect 38 -46 39 -44
rect 41 -46 43 -44
rect 38 -51 43 -46
rect 57 -35 70 -34
rect 57 -37 58 -35
rect 60 -37 62 -35
rect 64 -37 70 -35
rect 57 -38 70 -37
rect 57 -47 61 -38
rect 89 -42 93 -20
rect 88 -44 93 -42
rect 88 -46 89 -44
rect 91 -46 93 -44
rect 38 -53 39 -51
rect 41 -53 43 -51
rect 38 -55 43 -53
rect 88 -51 93 -46
rect 114 -11 136 -10
rect 114 -13 117 -11
rect 119 -13 136 -11
rect 114 -14 136 -13
rect 194 -11 199 -9
rect 194 -13 195 -11
rect 197 -13 199 -11
rect 114 -34 118 -14
rect 114 -36 120 -34
rect 114 -38 117 -36
rect 119 -38 120 -36
rect 114 -43 120 -38
rect 114 -45 117 -43
rect 119 -45 120 -43
rect 114 -47 120 -45
rect 147 -26 151 -17
rect 194 -15 199 -13
rect 138 -27 153 -26
rect 138 -29 139 -27
rect 141 -29 142 -27
rect 144 -29 149 -27
rect 151 -29 153 -27
rect 138 -30 153 -29
rect 163 -27 171 -25
rect 163 -29 168 -27
rect 170 -29 171 -27
rect 163 -31 171 -29
rect 163 -34 168 -31
rect 130 -35 168 -34
rect 130 -37 131 -35
rect 133 -37 168 -35
rect 130 -38 168 -37
rect 195 -37 199 -15
rect 194 -39 199 -37
rect 194 -41 195 -39
rect 197 -41 199 -39
rect 194 -46 199 -41
rect 194 -48 195 -46
rect 197 -48 199 -46
rect 194 -50 199 -48
rect 88 -53 89 -51
rect 91 -53 93 -51
rect 88 -55 93 -53
rect 186 -54 199 -50
rect -11 -64 203 -60
rect 3 -68 203 -64
<< alu2 >>
rect 38 61 134 62
rect 38 59 39 61
rect 41 59 131 61
rect 133 59 134 61
rect 38 58 134 59
rect 16 45 61 46
rect 16 43 17 45
rect 19 43 58 45
rect 60 43 61 45
rect 16 42 61 43
rect 130 45 134 46
rect 130 43 131 45
rect 133 43 134 45
rect 130 42 134 43
rect 14 28 18 29
rect 14 26 15 28
rect 17 26 18 28
rect 14 25 18 26
rect 64 28 68 29
rect 64 26 65 28
rect 67 26 68 28
rect 64 25 68 26
rect 147 28 151 29
rect 147 26 148 28
rect 150 26 151 28
rect 147 25 151 26
rect 132 21 136 22
rect 88 20 113 21
rect 88 18 89 20
rect 91 18 110 20
rect 112 18 113 20
rect 132 19 133 21
rect 135 19 136 21
rect 132 18 136 19
rect 88 17 113 18
rect 88 -10 151 -9
rect 88 -12 89 -10
rect 91 -12 148 -10
rect 150 -12 151 -10
rect 88 -13 151 -12
rect 14 -18 18 -17
rect 14 -20 15 -18
rect 17 -20 18 -18
rect 14 -21 18 -20
rect 64 -18 68 -17
rect 64 -20 65 -18
rect 67 -20 68 -18
rect 64 -21 68 -20
rect 132 -27 142 -26
rect 132 -29 133 -27
rect 135 -29 139 -27
rect 141 -29 142 -27
rect 132 -30 142 -29
rect 16 -35 61 -34
rect 16 -37 17 -35
rect 19 -37 58 -35
rect 60 -37 61 -35
rect 16 -38 61 -37
rect 109 -35 134 -34
rect 109 -37 110 -35
rect 112 -37 131 -35
rect 133 -37 134 -35
rect 109 -38 134 -37
<< alu3 >>
rect 130 61 134 62
rect 130 59 131 61
rect 133 59 134 61
rect 130 45 134 59
rect 130 43 131 45
rect 133 43 134 45
rect 130 42 134 43
rect 14 28 18 29
rect 14 26 15 28
rect 17 26 18 28
rect 14 -18 18 26
rect 14 -20 15 -18
rect 17 -20 18 -18
rect 14 -21 18 -20
rect 64 28 68 29
rect 64 26 65 28
rect 67 26 68 28
rect 64 -18 68 26
rect 147 28 151 29
rect 147 26 148 28
rect 150 26 151 28
rect 132 21 136 22
rect 64 -20 65 -18
rect 67 -20 68 -18
rect 64 -21 68 -20
rect 109 20 113 21
rect 109 18 110 20
rect 112 18 113 20
rect 109 -35 113 18
rect 132 19 133 21
rect 135 19 136 21
rect 132 -27 136 19
rect 147 -10 151 26
rect 147 -12 148 -10
rect 150 -12 151 -10
rect 147 -13 151 -12
rect 132 -29 133 -27
rect 135 -29 136 -27
rect 132 -30 136 -29
rect 109 -37 110 -35
rect 112 -37 113 -35
rect 109 -38 113 -37
<< nmos >>
rect 14 17 16 30
rect 21 17 23 30
rect 34 16 36 30
rect 64 17 66 30
rect 71 17 73 30
rect 84 16 86 30
rect 122 10 124 24
rect 133 10 135 30
rect 140 10 142 30
rect 160 16 162 30
rect 170 16 172 30
rect 180 13 182 23
rect 190 10 192 23
rect 14 -22 16 -9
rect 21 -22 23 -9
rect 34 -22 36 -8
rect 64 -22 66 -9
rect 71 -22 73 -9
rect 84 -22 86 -8
rect 122 -16 124 -2
rect 133 -22 135 -2
rect 140 -22 142 -2
rect 160 -22 162 -8
rect 170 -22 172 -8
rect 180 -15 182 -5
rect 190 -15 192 -2
<< pmos >>
rect 14 51 16 70
rect 24 51 26 70
rect 34 42 36 70
rect 64 51 66 70
rect 74 51 76 70
rect 84 42 86 70
rect 122 42 124 70
rect 132 42 134 70
rect 142 42 144 70
rect 160 42 162 67
rect 167 42 169 67
rect 177 45 179 58
rect 190 45 192 70
rect 14 -62 16 -43
rect 24 -62 26 -43
rect 34 -62 36 -34
rect 64 -62 66 -43
rect 74 -62 76 -43
rect 84 -62 86 -34
rect 122 -62 124 -34
rect 132 -62 134 -34
rect 142 -62 144 -34
rect 160 -59 162 -34
rect 167 -59 169 -34
rect 177 -50 179 -37
rect 190 -62 192 -37
<< polyct0 >>
rect 32 35 34 37
rect 82 35 84 37
rect 122 35 124 37
rect 132 35 134 37
rect 182 38 184 40
rect 188 28 190 30
rect 32 -29 34 -27
rect 82 -29 84 -27
rect 122 -29 124 -27
rect 132 -29 134 -27
rect 188 -22 190 -20
rect 182 -32 184 -30
<< polyct1 >>
rect 12 43 14 45
rect 62 43 64 45
rect 22 35 24 37
rect 72 35 74 37
rect 142 35 144 37
rect 149 35 151 37
rect 168 35 170 37
rect 22 -29 24 -27
rect 12 -37 14 -35
rect 72 -29 74 -27
rect 142 -29 144 -27
rect 149 -29 151 -27
rect 168 -29 170 -27
rect 62 -37 64 -35
<< ndifct0 >>
rect 9 19 11 21
rect 59 19 61 21
rect 128 12 130 14
rect 155 26 157 28
rect 145 19 147 21
rect 155 19 157 21
rect 165 26 167 28
rect 175 18 177 20
rect 185 15 187 17
rect 9 -13 11 -11
rect 59 -13 61 -11
rect 128 -6 130 -4
rect 145 -13 147 -11
rect 155 -13 157 -11
rect 155 -20 157 -18
rect 165 -20 167 -18
rect 175 -12 177 -10
rect 185 -9 187 -7
<< ndifct1 >>
rect 39 26 41 28
rect 39 18 41 20
rect 89 26 91 28
rect 89 18 91 20
rect 117 19 119 21
rect 28 9 30 11
rect 78 9 80 11
rect 195 19 197 21
rect 28 -3 30 -1
rect 78 -3 80 -1
rect 39 -12 41 -10
rect 39 -20 41 -18
rect 89 -12 91 -10
rect 117 -13 119 -11
rect 89 -20 91 -18
rect 195 -13 197 -11
<< pdifct0 >>
rect 9 66 11 68
rect 9 59 11 61
rect 19 60 21 62
rect 19 53 21 55
rect 29 66 31 68
rect 29 59 31 61
rect 59 66 61 68
rect 59 59 61 61
rect 69 60 71 62
rect 69 53 71 55
rect 79 66 81 68
rect 79 59 81 61
rect 127 66 129 68
rect 127 59 129 61
rect 137 58 139 60
rect 137 51 139 53
rect 149 66 151 68
rect 149 59 151 61
rect 184 66 186 68
rect 172 47 174 49
rect 9 -53 11 -51
rect 9 -60 11 -58
rect 19 -47 21 -45
rect 19 -54 21 -52
rect 29 -53 31 -51
rect 29 -60 31 -58
rect 59 -53 61 -51
rect 59 -60 61 -58
rect 69 -47 71 -45
rect 69 -54 71 -52
rect 79 -53 81 -51
rect 79 -60 81 -58
rect 127 -53 129 -51
rect 127 -60 129 -58
rect 137 -45 139 -43
rect 137 -52 139 -50
rect 149 -53 151 -51
rect 149 -60 151 -58
rect 172 -41 174 -39
rect 184 -60 186 -58
<< pdifct1 >>
rect 39 59 41 61
rect 39 52 41 54
rect 89 59 91 61
rect 89 52 91 54
rect 117 51 119 53
rect 117 44 119 46
rect 195 54 197 56
rect 195 47 197 49
rect 39 -46 41 -44
rect 39 -53 41 -51
rect 117 -38 119 -36
rect 89 -46 91 -44
rect 117 -45 119 -43
rect 89 -53 91 -51
rect 195 -41 197 -39
rect 195 -48 197 -46
<< alu0 >>
rect 7 66 9 68
rect 11 66 13 68
rect 7 61 13 66
rect 27 66 29 68
rect 31 66 33 68
rect 7 59 9 61
rect 11 59 13 61
rect 7 58 13 59
rect 17 62 23 63
rect 17 60 19 62
rect 21 60 23 62
rect 17 55 23 60
rect 27 61 33 66
rect 57 66 59 68
rect 61 66 63 68
rect 27 59 29 61
rect 31 59 33 61
rect 27 58 33 59
rect 17 53 19 55
rect 21 54 23 55
rect 57 61 63 66
rect 77 66 79 68
rect 81 66 83 68
rect 57 59 59 61
rect 61 59 63 61
rect 57 58 63 59
rect 67 62 73 63
rect 67 60 69 62
rect 71 60 73 62
rect 67 55 73 60
rect 77 61 83 66
rect 125 66 127 68
rect 129 66 131 68
rect 77 59 79 61
rect 81 59 83 61
rect 77 58 83 59
rect 21 53 31 54
rect 17 50 31 53
rect 27 46 31 50
rect 27 42 35 46
rect 31 37 35 42
rect 31 35 32 37
rect 34 35 35 37
rect 31 30 35 35
rect 23 26 35 30
rect 23 22 27 26
rect 38 23 39 30
rect 67 53 69 55
rect 71 54 73 55
rect 125 61 131 66
rect 147 66 149 68
rect 151 66 153 68
rect 125 59 127 61
rect 129 59 131 61
rect 125 58 131 59
rect 136 60 140 62
rect 136 58 137 60
rect 139 58 140 60
rect 147 61 153 66
rect 182 66 184 68
rect 186 66 188 68
rect 182 65 188 66
rect 147 59 149 61
rect 151 59 153 61
rect 147 58 153 59
rect 71 53 81 54
rect 67 50 81 53
rect 77 46 81 50
rect 77 42 85 46
rect 81 37 85 42
rect 81 35 82 37
rect 84 35 85 37
rect 81 30 85 35
rect 73 26 85 30
rect 7 21 27 22
rect 7 19 9 21
rect 11 19 27 21
rect 7 18 27 19
rect 73 22 77 26
rect 88 23 89 30
rect 57 21 77 22
rect 57 19 59 21
rect 61 19 77 21
rect 57 18 77 19
rect 136 54 140 58
rect 159 54 183 58
rect 123 53 163 54
rect 123 51 137 53
rect 139 51 163 53
rect 123 50 163 51
rect 123 39 127 50
rect 171 49 175 51
rect 179 50 185 54
rect 171 47 172 49
rect 174 47 175 49
rect 171 46 175 47
rect 171 42 178 46
rect 121 37 127 39
rect 121 35 122 37
rect 124 35 127 37
rect 121 33 127 35
rect 131 37 135 42
rect 131 35 132 37
rect 134 35 135 37
rect 131 33 135 35
rect 123 30 127 33
rect 123 26 143 30
rect 139 22 143 26
rect 174 31 178 42
rect 181 40 185 50
rect 181 38 182 40
rect 184 38 185 40
rect 181 36 185 38
rect 174 30 192 31
rect 154 28 158 30
rect 174 29 188 30
rect 154 26 155 28
rect 157 26 158 28
rect 139 21 149 22
rect 139 19 145 21
rect 147 19 149 21
rect 139 18 149 19
rect 154 21 158 26
rect 163 28 188 29
rect 190 28 192 30
rect 163 26 165 28
rect 167 27 192 28
rect 167 26 178 27
rect 163 25 178 26
rect 154 19 155 21
rect 157 20 179 21
rect 157 19 175 20
rect 154 18 175 19
rect 177 18 179 20
rect 154 17 179 18
rect 184 17 188 19
rect 184 15 185 17
rect 187 15 188 17
rect 126 14 132 15
rect 126 12 128 14
rect 130 12 132 14
rect 184 12 188 15
rect 126 -6 128 -4
rect 130 -6 132 -4
rect 126 -7 132 -6
rect 184 -7 188 -4
rect 184 -9 185 -7
rect 187 -9 188 -7
rect 154 -10 179 -9
rect 7 -11 27 -10
rect 7 -13 9 -11
rect 11 -13 27 -11
rect 7 -14 27 -13
rect 23 -18 27 -14
rect 57 -11 77 -10
rect 57 -13 59 -11
rect 61 -13 77 -11
rect 57 -14 77 -13
rect 23 -22 35 -18
rect 38 -22 39 -15
rect 31 -27 35 -22
rect 31 -29 32 -27
rect 34 -29 35 -27
rect 31 -34 35 -29
rect 27 -38 35 -34
rect 27 -42 31 -38
rect 73 -18 77 -14
rect 73 -22 85 -18
rect 88 -22 89 -15
rect 81 -27 85 -22
rect 81 -29 82 -27
rect 84 -29 85 -27
rect 81 -34 85 -29
rect 17 -45 31 -42
rect 17 -47 19 -45
rect 21 -46 31 -45
rect 21 -47 23 -46
rect 7 -51 13 -50
rect 7 -53 9 -51
rect 11 -53 13 -51
rect 7 -58 13 -53
rect 17 -52 23 -47
rect 17 -54 19 -52
rect 21 -54 23 -52
rect 17 -55 23 -54
rect 27 -51 33 -50
rect 27 -53 29 -51
rect 31 -53 33 -51
rect 7 -60 9 -58
rect 11 -60 13 -58
rect 27 -58 33 -53
rect 77 -38 85 -34
rect 77 -42 81 -38
rect 67 -45 81 -42
rect 67 -47 69 -45
rect 71 -46 81 -45
rect 71 -47 73 -46
rect 57 -51 63 -50
rect 57 -53 59 -51
rect 61 -53 63 -51
rect 27 -60 29 -58
rect 31 -60 33 -58
rect 57 -58 63 -53
rect 67 -52 73 -47
rect 67 -54 69 -52
rect 71 -54 73 -52
rect 67 -55 73 -54
rect 77 -51 83 -50
rect 77 -53 79 -51
rect 81 -53 83 -51
rect 57 -60 59 -58
rect 61 -60 63 -58
rect 77 -58 83 -53
rect 139 -11 149 -10
rect 139 -13 145 -11
rect 147 -13 149 -11
rect 139 -14 149 -13
rect 154 -11 175 -10
rect 154 -13 155 -11
rect 157 -12 175 -11
rect 177 -12 179 -10
rect 184 -11 188 -9
rect 157 -13 179 -12
rect 139 -18 143 -14
rect 123 -22 143 -18
rect 123 -25 127 -22
rect 121 -27 127 -25
rect 121 -29 122 -27
rect 124 -29 127 -27
rect 121 -31 127 -29
rect 123 -42 127 -31
rect 131 -27 135 -25
rect 154 -18 158 -13
rect 154 -20 155 -18
rect 157 -20 158 -18
rect 154 -22 158 -20
rect 163 -18 178 -17
rect 163 -20 165 -18
rect 167 -19 178 -18
rect 167 -20 192 -19
rect 163 -21 188 -20
rect 174 -22 188 -21
rect 190 -22 192 -20
rect 174 -23 192 -22
rect 131 -29 132 -27
rect 134 -29 135 -27
rect 131 -34 135 -29
rect 174 -34 178 -23
rect 171 -38 178 -34
rect 181 -30 185 -28
rect 181 -32 182 -30
rect 184 -32 185 -30
rect 171 -39 175 -38
rect 171 -41 172 -39
rect 174 -41 175 -39
rect 123 -43 163 -42
rect 171 -43 175 -41
rect 181 -42 185 -32
rect 123 -45 137 -43
rect 139 -45 163 -43
rect 123 -46 163 -45
rect 179 -46 185 -42
rect 136 -50 140 -46
rect 159 -50 183 -46
rect 125 -51 131 -50
rect 125 -53 127 -51
rect 129 -53 131 -51
rect 77 -60 79 -58
rect 81 -60 83 -58
rect 125 -58 131 -53
rect 136 -52 137 -50
rect 139 -52 140 -50
rect 136 -54 140 -52
rect 147 -51 153 -50
rect 147 -53 149 -51
rect 151 -53 153 -51
rect 125 -60 127 -58
rect 129 -60 131 -58
rect 147 -58 153 -53
rect 147 -60 149 -58
rect 151 -60 153 -58
rect 182 -58 188 -57
rect 182 -60 184 -58
rect 186 -60 188 -58
<< via1 >>
rect 39 59 41 61
rect 17 43 19 45
rect 15 26 17 28
rect 58 43 60 45
rect 65 26 67 28
rect 89 18 91 20
rect 131 43 133 45
rect 148 26 150 28
rect 133 19 135 21
rect 15 -20 17 -18
rect 17 -37 19 -35
rect 65 -20 67 -18
rect 89 -12 91 -10
rect 58 -37 60 -35
rect 139 -29 141 -27
rect 131 -37 133 -35
<< via2 >>
rect 131 59 133 61
rect 131 43 133 45
rect 15 26 17 28
rect 65 26 67 28
rect 148 26 150 28
rect 110 18 112 20
rect 133 19 135 21
rect 148 -12 150 -10
rect 15 -20 17 -18
rect 65 -20 67 -18
rect 133 -29 135 -27
rect 110 -37 112 -35
<< labels >>
rlabel alu1 25 8 25 8 4 vss
rlabel alu1 25 72 25 72 4 vdd
rlabel alu1 25 0 25 0 2 vss
rlabel alu0 20 -48 20 -48 2 zn
rlabel alu0 17 -12 17 -12 2 zn
rlabel polyct0 33 -28 33 -28 2 zn
rlabel alu1 75 8 75 8 4 vss
rlabel alu1 75 72 75 72 4 vdd
rlabel alu1 75 0 75 0 2 vss
rlabel alu1 153 0 153 0 2 vss
rlabel alu0 183 45 183 45 4 con
rlabel alu0 171 27 171 27 4 son
rlabel alu0 183 29 183 29 4 son
rlabel alu0 173 46 173 46 4 son
rlabel alu0 167 19 167 19 4 n2
rlabel alu0 144 20 144 20 4 con
rlabel alu0 156 23 156 23 4 n2
rlabel alu0 125 40 125 40 4 con
rlabel alu0 143 52 143 52 4 con
rlabel alu0 138 56 138 56 4 con
rlabel alu1 153 8 153 8 4 vss
rlabel alu1 133 20 133 20 4 co
rlabel alu1 153 72 153 72 4 vdd
rlabel alu1 117 20 117 20 4 co
rlabel alu1 125 20 125 20 4 co
rlabel alu1 117 48 117 48 4 co
rlabel alu1 17 -24 17 -24 1 a2
rlabel alu1 25 -28 25 -28 1 a2
rlabel alu1 17 -36 17 -36 1 b2
rlabel alu1 9 -44 9 -44 1 b2
rlabel alu1 17 32 17 32 1 a2
rlabel alu1 25 36 25 36 1 a2
rlabel alu1 17 44 17 44 1 b3
rlabel alu1 9 52 9 52 1 b3
rlabel alu1 59 52 59 52 1 b3
rlabel alu1 67 44 67 44 1 b3
rlabel alu1 67 32 67 32 1 a3
rlabel alu1 75 36 75 36 1 a3
rlabel alu1 59 -44 59 -44 1 b2
rlabel alu1 67 -36 67 -36 1 b2
rlabel alu1 75 -28 75 -28 1 a3
rlabel alu1 41 40 41 40 1 z2
rlabel alu1 91 40 91 40 1 z1
rlabel alu1 91 -32 91 -32 1 z3
rlabel alu1 33 20 33 20 1 z2
rlabel alu1 83 20 83 20 1 z1
rlabel alu1 83 -12 83 -12 1 z3
rlabel alu1 197 36 197 36 1 p1
rlabel alu1 189 60 189 60 1 p1
rlabel alu1 33 -12 33 -12 1 p0
rlabel alu1 41 -32 41 -32 1 p0
rlabel alu1 197 -28 197 -28 1 p2
rlabel alu1 189 -52 189 -52 1 p2
rlabel polyct0 83 -28 83 -28 2 zn_uq0
rlabel alu0 67 -12 67 -12 2 zn_uq0
rlabel alu0 70 -48 70 -48 2 zn_uq0
rlabel alu0 70 56 70 56 4 zn_uq1
rlabel alu0 67 20 67 20 4 zn_uq1
rlabel polyct0 83 36 83 36 4 zn_uq1
rlabel alu0 20 56 20 56 4 zn_uq2
rlabel alu0 17 20 17 20 4 zn_uq2
rlabel polyct0 33 36 33 36 4 zn_uq2
rlabel alu0 167 -11 167 -11 2 n2_uq0
rlabel alu0 156 -15 156 -15 2 n2_uq0
rlabel alu0 171 -19 171 -19 2 son_uq0
rlabel alu0 183 -21 183 -21 2 son_uq0
rlabel alu0 173 -38 173 -38 2 son_uq0
rlabel alu0 183 -37 183 -37 2 con_uq0
rlabel alu0 144 -12 144 -12 2 con_uq0
rlabel alu0 125 -32 125 -32 2 con_uq0
rlabel alu0 143 -44 143 -44 2 con_uq0
rlabel alu0 138 -48 138 -48 2 con_uq0
rlabel nmos 66 -22 66 -22 1 a3_uq0
rlabel alu1 75 -28 75 -28 1 a2_uq0
rlabel alu1 117 -40 117 -40 1 p3
rlabel alu1 116 -29 116 -29 1 p3
<< end >>
